VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO multiply_4
  CLASS BLOCK ;
  FOREIGN multiply_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 998.810 BY 1000.125 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.920 0.000 499.200 4.000 ;
    END
  END clk
  PIN m_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.740 996.000 1.020 1000.000 ;
    END
  END m_in[0]
  PIN m_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.680 996.000 386.960 1000.000 ;
    END
  END m_in[100]
  PIN m_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.360 996.000 390.640 1000.000 ;
    END
  END m_in[101]
  PIN m_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.500 996.000 394.780 1000.000 ;
    END
  END m_in[102]
  PIN m_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.180 996.000 398.460 1000.000 ;
    END
  END m_in[103]
  PIN m_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.860 996.000 402.140 1000.000 ;
    END
  END m_in[104]
  PIN m_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.000 996.000 406.280 1000.000 ;
    END
  END m_in[105]
  PIN m_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.680 996.000 409.960 1000.000 ;
    END
  END m_in[106]
  PIN m_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.820 996.000 414.100 1000.000 ;
    END
  END m_in[107]
  PIN m_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.500 996.000 417.780 1000.000 ;
    END
  END m_in[108]
  PIN m_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.180 996.000 421.460 1000.000 ;
    END
  END m_in[109]
  PIN m_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.920 996.000 39.200 1000.000 ;
    END
  END m_in[10]
  PIN m_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.320 996.000 425.600 1000.000 ;
    END
  END m_in[110]
  PIN m_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.000 996.000 429.280 1000.000 ;
    END
  END m_in[111]
  PIN m_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.140 996.000 433.420 1000.000 ;
    END
  END m_in[112]
  PIN m_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.820 996.000 437.100 1000.000 ;
    END
  END m_in[113]
  PIN m_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.500 996.000 440.780 1000.000 ;
    END
  END m_in[114]
  PIN m_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.640 996.000 444.920 1000.000 ;
    END
  END m_in[115]
  PIN m_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.320 996.000 448.600 1000.000 ;
    END
  END m_in[116]
  PIN m_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.460 996.000 452.740 1000.000 ;
    END
  END m_in[117]
  PIN m_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.140 996.000 456.420 1000.000 ;
    END
  END m_in[118]
  PIN m_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.820 996.000 460.100 1000.000 ;
    END
  END m_in[119]
  PIN m_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.060 996.000 43.340 1000.000 ;
    END
  END m_in[11]
  PIN m_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.960 996.000 464.240 1000.000 ;
    END
  END m_in[120]
  PIN m_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.640 996.000 467.920 1000.000 ;
    END
  END m_in[121]
  PIN m_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.780 996.000 472.060 1000.000 ;
    END
  END m_in[122]
  PIN m_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.460 996.000 475.740 1000.000 ;
    END
  END m_in[123]
  PIN m_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.140 996.000 479.420 1000.000 ;
    END
  END m_in[124]
  PIN m_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.280 996.000 483.560 1000.000 ;
    END
  END m_in[125]
  PIN m_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.960 996.000 487.240 1000.000 ;
    END
  END m_in[126]
  PIN m_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.100 996.000 491.380 1000.000 ;
    END
  END m_in[127]
  PIN m_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.780 996.000 495.060 1000.000 ;
    END
  END m_in[128]
  PIN m_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.460 996.000 498.740 1000.000 ;
    END
  END m_in[129]
  PIN m_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.740 996.000 47.020 1000.000 ;
    END
  END m_in[12]
  PIN m_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.600 996.000 502.880 1000.000 ;
    END
  END m_in[130]
  PIN m_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.280 996.000 506.560 1000.000 ;
    END
  END m_in[131]
  PIN m_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.960 996.000 510.240 1000.000 ;
    END
  END m_in[132]
  PIN m_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.100 996.000 514.380 1000.000 ;
    END
  END m_in[133]
  PIN m_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.780 996.000 518.060 1000.000 ;
    END
  END m_in[134]
  PIN m_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.920 996.000 522.200 1000.000 ;
    END
  END m_in[135]
  PIN m_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.600 996.000 525.880 1000.000 ;
    END
  END m_in[136]
  PIN m_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.280 996.000 529.560 1000.000 ;
    END
  END m_in[137]
  PIN m_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.420 996.000 533.700 1000.000 ;
    END
  END m_in[138]
  PIN m_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.100 996.000 537.380 1000.000 ;
    END
  END m_in[139]
  PIN m_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.880 996.000 51.160 1000.000 ;
    END
  END m_in[13]
  PIN m_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.240 996.000 541.520 1000.000 ;
    END
  END m_in[140]
  PIN m_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.920 996.000 545.200 1000.000 ;
    END
  END m_in[141]
  PIN m_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.600 996.000 548.880 1000.000 ;
    END
  END m_in[142]
  PIN m_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.740 996.000 553.020 1000.000 ;
    END
  END m_in[143]
  PIN m_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.420 996.000 556.700 1000.000 ;
    END
  END m_in[144]
  PIN m_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.560 996.000 560.840 1000.000 ;
    END
  END m_in[145]
  PIN m_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.240 996.000 564.520 1000.000 ;
    END
  END m_in[146]
  PIN m_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.920 996.000 568.200 1000.000 ;
    END
  END m_in[147]
  PIN m_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.060 996.000 572.340 1000.000 ;
    END
  END m_in[148]
  PIN m_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.740 996.000 576.020 1000.000 ;
    END
  END m_in[149]
  PIN m_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.560 996.000 54.840 1000.000 ;
    END
  END m_in[14]
  PIN m_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.880 996.000 580.160 1000.000 ;
    END
  END m_in[150]
  PIN m_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.560 996.000 583.840 1000.000 ;
    END
  END m_in[151]
  PIN m_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.240 996.000 587.520 1000.000 ;
    END
  END m_in[152]
  PIN m_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.380 996.000 591.660 1000.000 ;
    END
  END m_in[153]
  PIN m_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.060 996.000 595.340 1000.000 ;
    END
  END m_in[154]
  PIN m_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.200 996.000 599.480 1000.000 ;
    END
  END m_in[155]
  PIN m_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.880 996.000 603.160 1000.000 ;
    END
  END m_in[156]
  PIN m_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.560 996.000 606.840 1000.000 ;
    END
  END m_in[157]
  PIN m_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.700 996.000 610.980 1000.000 ;
    END
  END m_in[158]
  PIN m_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.380 996.000 614.660 1000.000 ;
    END
  END m_in[159]
  PIN m_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.240 996.000 58.520 1000.000 ;
    END
  END m_in[15]
  PIN m_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.520 996.000 618.800 1000.000 ;
    END
  END m_in[160]
  PIN m_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.200 996.000 622.480 1000.000 ;
    END
  END m_in[161]
  PIN m_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.880 996.000 626.160 1000.000 ;
    END
  END m_in[162]
  PIN m_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.020 996.000 630.300 1000.000 ;
    END
  END m_in[163]
  PIN m_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.700 996.000 633.980 1000.000 ;
    END
  END m_in[164]
  PIN m_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.380 996.000 637.660 1000.000 ;
    END
  END m_in[165]
  PIN m_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.520 996.000 641.800 1000.000 ;
    END
  END m_in[166]
  PIN m_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.200 996.000 645.480 1000.000 ;
    END
  END m_in[167]
  PIN m_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.340 996.000 649.620 1000.000 ;
    END
  END m_in[168]
  PIN m_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.020 996.000 653.300 1000.000 ;
    END
  END m_in[169]
  PIN m_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.380 996.000 62.660 1000.000 ;
    END
  END m_in[16]
  PIN m_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.700 996.000 656.980 1000.000 ;
    END
  END m_in[170]
  PIN m_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.840 996.000 661.120 1000.000 ;
    END
  END m_in[171]
  PIN m_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.520 996.000 664.800 1000.000 ;
    END
  END m_in[172]
  PIN m_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.660 996.000 668.940 1000.000 ;
    END
  END m_in[173]
  PIN m_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.340 996.000 672.620 1000.000 ;
    END
  END m_in[174]
  PIN m_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.020 996.000 676.300 1000.000 ;
    END
  END m_in[175]
  PIN m_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.160 996.000 680.440 1000.000 ;
    END
  END m_in[176]
  PIN m_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.840 996.000 684.120 1000.000 ;
    END
  END m_in[177]
  PIN m_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.980 996.000 688.260 1000.000 ;
    END
  END m_in[178]
  PIN m_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.660 996.000 691.940 1000.000 ;
    END
  END m_in[179]
  PIN m_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.060 996.000 66.340 1000.000 ;
    END
  END m_in[17]
  PIN m_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.340 996.000 695.620 1000.000 ;
    END
  END m_in[180]
  PIN m_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.480 996.000 699.760 1000.000 ;
    END
  END m_in[181]
  PIN m_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.160 996.000 703.440 1000.000 ;
    END
  END m_in[182]
  PIN m_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.300 996.000 707.580 1000.000 ;
    END
  END m_in[183]
  PIN m_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.980 996.000 711.260 1000.000 ;
    END
  END m_in[184]
  PIN m_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.660 996.000 714.940 1000.000 ;
    END
  END m_in[185]
  PIN m_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.800 996.000 719.080 1000.000 ;
    END
  END m_in[186]
  PIN m_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.480 996.000 722.760 1000.000 ;
    END
  END m_in[187]
  PIN m_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.620 996.000 726.900 1000.000 ;
    END
  END m_in[188]
  PIN m_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.300 996.000 730.580 1000.000 ;
    END
  END m_in[189]
  PIN m_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.200 996.000 70.480 1000.000 ;
    END
  END m_in[18]
  PIN m_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.980 996.000 734.260 1000.000 ;
    END
  END m_in[190]
  PIN m_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.120 996.000 738.400 1000.000 ;
    END
  END m_in[191]
  PIN m_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.800 996.000 742.080 1000.000 ;
    END
  END m_in[192]
  PIN m_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.940 996.000 746.220 1000.000 ;
    END
  END m_in[193]
  PIN m_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.620 996.000 749.900 1000.000 ;
    END
  END m_in[194]
  PIN m_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.300 996.000 753.580 1000.000 ;
    END
  END m_in[195]
  PIN m_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.440 996.000 757.720 1000.000 ;
    END
  END m_in[196]
  PIN m_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.120 996.000 761.400 1000.000 ;
    END
  END m_in[197]
  PIN m_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.800 996.000 765.080 1000.000 ;
    END
  END m_in[198]
  PIN m_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.940 996.000 769.220 1000.000 ;
    END
  END m_in[199]
  PIN m_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.880 996.000 74.160 1000.000 ;
    END
  END m_in[19]
  PIN m_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.420 996.000 4.700 1000.000 ;
    END
  END m_in[1]
  PIN m_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.620 996.000 772.900 1000.000 ;
    END
  END m_in[200]
  PIN m_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.760 996.000 777.040 1000.000 ;
    END
  END m_in[201]
  PIN m_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.440 996.000 780.720 1000.000 ;
    END
  END m_in[202]
  PIN m_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.120 996.000 784.400 1000.000 ;
    END
  END m_in[203]
  PIN m_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.260 996.000 788.540 1000.000 ;
    END
  END m_in[204]
  PIN m_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.940 996.000 792.220 1000.000 ;
    END
  END m_in[205]
  PIN m_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.080 996.000 796.360 1000.000 ;
    END
  END m_in[206]
  PIN m_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.760 996.000 800.040 1000.000 ;
    END
  END m_in[207]
  PIN m_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.440 996.000 803.720 1000.000 ;
    END
  END m_in[208]
  PIN m_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.580 996.000 807.860 1000.000 ;
    END
  END m_in[209]
  PIN m_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.560 996.000 77.840 1000.000 ;
    END
  END m_in[20]
  PIN m_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.260 996.000 811.540 1000.000 ;
    END
  END m_in[210]
  PIN m_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.400 996.000 815.680 1000.000 ;
    END
  END m_in[211]
  PIN m_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.080 996.000 819.360 1000.000 ;
    END
  END m_in[212]
  PIN m_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.760 996.000 823.040 1000.000 ;
    END
  END m_in[213]
  PIN m_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.900 996.000 827.180 1000.000 ;
    END
  END m_in[214]
  PIN m_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.580 996.000 830.860 1000.000 ;
    END
  END m_in[215]
  PIN m_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.720 996.000 835.000 1000.000 ;
    END
  END m_in[216]
  PIN m_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.400 996.000 838.680 1000.000 ;
    END
  END m_in[217]
  PIN m_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.080 996.000 842.360 1000.000 ;
    END
  END m_in[218]
  PIN m_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.220 996.000 846.500 1000.000 ;
    END
  END m_in[219]
  PIN m_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.700 996.000 81.980 1000.000 ;
    END
  END m_in[21]
  PIN m_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.900 996.000 850.180 1000.000 ;
    END
  END m_in[220]
  PIN m_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.040 996.000 854.320 1000.000 ;
    END
  END m_in[221]
  PIN m_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.720 996.000 858.000 1000.000 ;
    END
  END m_in[222]
  PIN m_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.400 996.000 861.680 1000.000 ;
    END
  END m_in[223]
  PIN m_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.540 996.000 865.820 1000.000 ;
    END
  END m_in[224]
  PIN m_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.220 996.000 869.500 1000.000 ;
    END
  END m_in[225]
  PIN m_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.360 996.000 873.640 1000.000 ;
    END
  END m_in[226]
  PIN m_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.040 996.000 877.320 1000.000 ;
    END
  END m_in[227]
  PIN m_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.720 996.000 881.000 1000.000 ;
    END
  END m_in[228]
  PIN m_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.860 996.000 885.140 1000.000 ;
    END
  END m_in[229]
  PIN m_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.380 996.000 85.660 1000.000 ;
    END
  END m_in[22]
  PIN m_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.540 996.000 888.820 1000.000 ;
    END
  END m_in[230]
  PIN m_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.220 996.000 892.500 1000.000 ;
    END
  END m_in[231]
  PIN m_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.360 996.000 896.640 1000.000 ;
    END
  END m_in[232]
  PIN m_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.040 996.000 900.320 1000.000 ;
    END
  END m_in[233]
  PIN m_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.180 996.000 904.460 1000.000 ;
    END
  END m_in[234]
  PIN m_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.860 996.000 908.140 1000.000 ;
    END
  END m_in[235]
  PIN m_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.540 996.000 911.820 1000.000 ;
    END
  END m_in[236]
  PIN m_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.680 996.000 915.960 1000.000 ;
    END
  END m_in[237]
  PIN m_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.360 996.000 919.640 1000.000 ;
    END
  END m_in[238]
  PIN m_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.500 996.000 923.780 1000.000 ;
    END
  END m_in[239]
  PIN m_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.520 996.000 89.800 1000.000 ;
    END
  END m_in[23]
  PIN m_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.180 996.000 927.460 1000.000 ;
    END
  END m_in[240]
  PIN m_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.860 996.000 931.140 1000.000 ;
    END
  END m_in[241]
  PIN m_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.000 996.000 935.280 1000.000 ;
    END
  END m_in[242]
  PIN m_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.680 996.000 938.960 1000.000 ;
    END
  END m_in[243]
  PIN m_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.820 996.000 943.100 1000.000 ;
    END
  END m_in[244]
  PIN m_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.500 996.000 946.780 1000.000 ;
    END
  END m_in[245]
  PIN m_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.180 996.000 950.460 1000.000 ;
    END
  END m_in[246]
  PIN m_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.320 996.000 954.600 1000.000 ;
    END
  END m_in[247]
  PIN m_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.000 996.000 958.280 1000.000 ;
    END
  END m_in[248]
  PIN m_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.140 996.000 962.420 1000.000 ;
    END
  END m_in[249]
  PIN m_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.200 996.000 93.480 1000.000 ;
    END
  END m_in[24]
  PIN m_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.820 996.000 966.100 1000.000 ;
    END
  END m_in[250]
  PIN m_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.500 996.000 969.780 1000.000 ;
    END
  END m_in[251]
  PIN m_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 973.640 996.000 973.920 1000.000 ;
    END
  END m_in[252]
  PIN m_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.320 996.000 977.600 1000.000 ;
    END
  END m_in[253]
  PIN m_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.460 996.000 981.740 1000.000 ;
    END
  END m_in[254]
  PIN m_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.140 996.000 985.420 1000.000 ;
    END
  END m_in[255]
  PIN m_in[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.820 996.000 989.100 1000.000 ;
    END
  END m_in[256]
  PIN m_in[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.960 996.000 993.240 1000.000 ;
    END
  END m_in[257]
  PIN m_in[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.640 996.000 996.920 1000.000 ;
    END
  END m_in[258]
  PIN m_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.880 996.000 97.160 1000.000 ;
    END
  END m_in[25]
  PIN m_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.020 996.000 101.300 1000.000 ;
    END
  END m_in[26]
  PIN m_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.700 996.000 104.980 1000.000 ;
    END
  END m_in[27]
  PIN m_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.840 996.000 109.120 1000.000 ;
    END
  END m_in[28]
  PIN m_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.520 996.000 112.800 1000.000 ;
    END
  END m_in[29]
  PIN m_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.100 996.000 8.380 1000.000 ;
    END
  END m_in[2]
  PIN m_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.200 996.000 116.480 1000.000 ;
    END
  END m_in[30]
  PIN m_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.340 996.000 120.620 1000.000 ;
    END
  END m_in[31]
  PIN m_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.020 996.000 124.300 1000.000 ;
    END
  END m_in[32]
  PIN m_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.700 996.000 127.980 1000.000 ;
    END
  END m_in[33]
  PIN m_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.840 996.000 132.120 1000.000 ;
    END
  END m_in[34]
  PIN m_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.520 996.000 135.800 1000.000 ;
    END
  END m_in[35]
  PIN m_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.660 996.000 139.940 1000.000 ;
    END
  END m_in[36]
  PIN m_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.340 996.000 143.620 1000.000 ;
    END
  END m_in[37]
  PIN m_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.020 996.000 147.300 1000.000 ;
    END
  END m_in[38]
  PIN m_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.160 996.000 151.440 1000.000 ;
    END
  END m_in[39]
  PIN m_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.240 996.000 12.520 1000.000 ;
    END
  END m_in[3]
  PIN m_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.840 996.000 155.120 1000.000 ;
    END
  END m_in[40]
  PIN m_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.980 996.000 159.260 1000.000 ;
    END
  END m_in[41]
  PIN m_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.660 996.000 162.940 1000.000 ;
    END
  END m_in[42]
  PIN m_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.340 996.000 166.620 1000.000 ;
    END
  END m_in[43]
  PIN m_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.480 996.000 170.760 1000.000 ;
    END
  END m_in[44]
  PIN m_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.160 996.000 174.440 1000.000 ;
    END
  END m_in[45]
  PIN m_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.300 996.000 178.580 1000.000 ;
    END
  END m_in[46]
  PIN m_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.980 996.000 182.260 1000.000 ;
    END
  END m_in[47]
  PIN m_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.660 996.000 185.940 1000.000 ;
    END
  END m_in[48]
  PIN m_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.800 996.000 190.080 1000.000 ;
    END
  END m_in[49]
  PIN m_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.920 996.000 16.200 1000.000 ;
    END
  END m_in[4]
  PIN m_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.480 996.000 193.760 1000.000 ;
    END
  END m_in[50]
  PIN m_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.620 996.000 197.900 1000.000 ;
    END
  END m_in[51]
  PIN m_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.300 996.000 201.580 1000.000 ;
    END
  END m_in[52]
  PIN m_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.980 996.000 205.260 1000.000 ;
    END
  END m_in[53]
  PIN m_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.120 996.000 209.400 1000.000 ;
    END
  END m_in[54]
  PIN m_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.800 996.000 213.080 1000.000 ;
    END
  END m_in[55]
  PIN m_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.940 996.000 217.220 1000.000 ;
    END
  END m_in[56]
  PIN m_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.620 996.000 220.900 1000.000 ;
    END
  END m_in[57]
  PIN m_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.300 996.000 224.580 1000.000 ;
    END
  END m_in[58]
  PIN m_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.440 996.000 228.720 1000.000 ;
    END
  END m_in[59]
  PIN m_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.600 996.000 19.880 1000.000 ;
    END
  END m_in[5]
  PIN m_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.120 996.000 232.400 1000.000 ;
    END
  END m_in[60]
  PIN m_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.260 996.000 236.540 1000.000 ;
    END
  END m_in[61]
  PIN m_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.940 996.000 240.220 1000.000 ;
    END
  END m_in[62]
  PIN m_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.620 996.000 243.900 1000.000 ;
    END
  END m_in[63]
  PIN m_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.760 996.000 248.040 1000.000 ;
    END
  END m_in[64]
  PIN m_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.440 996.000 251.720 1000.000 ;
    END
  END m_in[65]
  PIN m_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.120 996.000 255.400 1000.000 ;
    END
  END m_in[66]
  PIN m_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.260 996.000 259.540 1000.000 ;
    END
  END m_in[67]
  PIN m_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.940 996.000 263.220 1000.000 ;
    END
  END m_in[68]
  PIN m_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.080 996.000 267.360 1000.000 ;
    END
  END m_in[69]
  PIN m_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.740 996.000 24.020 1000.000 ;
    END
  END m_in[6]
  PIN m_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.760 996.000 271.040 1000.000 ;
    END
  END m_in[70]
  PIN m_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.440 996.000 274.720 1000.000 ;
    END
  END m_in[71]
  PIN m_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.580 996.000 278.860 1000.000 ;
    END
  END m_in[72]
  PIN m_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.260 996.000 282.540 1000.000 ;
    END
  END m_in[73]
  PIN m_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.400 996.000 286.680 1000.000 ;
    END
  END m_in[74]
  PIN m_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.080 996.000 290.360 1000.000 ;
    END
  END m_in[75]
  PIN m_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.760 996.000 294.040 1000.000 ;
    END
  END m_in[76]
  PIN m_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.900 996.000 298.180 1000.000 ;
    END
  END m_in[77]
  PIN m_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.580 996.000 301.860 1000.000 ;
    END
  END m_in[78]
  PIN m_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.720 996.000 306.000 1000.000 ;
    END
  END m_in[79]
  PIN m_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.420 996.000 27.700 1000.000 ;
    END
  END m_in[7]
  PIN m_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.400 996.000 309.680 1000.000 ;
    END
  END m_in[80]
  PIN m_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.080 996.000 313.360 1000.000 ;
    END
  END m_in[81]
  PIN m_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.220 996.000 317.500 1000.000 ;
    END
  END m_in[82]
  PIN m_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.900 996.000 321.180 1000.000 ;
    END
  END m_in[83]
  PIN m_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.040 996.000 325.320 1000.000 ;
    END
  END m_in[84]
  PIN m_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.720 996.000 329.000 1000.000 ;
    END
  END m_in[85]
  PIN m_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.400 996.000 332.680 1000.000 ;
    END
  END m_in[86]
  PIN m_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.540 996.000 336.820 1000.000 ;
    END
  END m_in[87]
  PIN m_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.220 996.000 340.500 1000.000 ;
    END
  END m_in[88]
  PIN m_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.360 996.000 344.640 1000.000 ;
    END
  END m_in[89]
  PIN m_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.560 996.000 31.840 1000.000 ;
    END
  END m_in[8]
  PIN m_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.040 996.000 348.320 1000.000 ;
    END
  END m_in[90]
  PIN m_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.720 996.000 352.000 1000.000 ;
    END
  END m_in[91]
  PIN m_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.860 996.000 356.140 1000.000 ;
    END
  END m_in[92]
  PIN m_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.540 996.000 359.820 1000.000 ;
    END
  END m_in[93]
  PIN m_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.680 996.000 363.960 1000.000 ;
    END
  END m_in[94]
  PIN m_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.360 996.000 367.640 1000.000 ;
    END
  END m_in[95]
  PIN m_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.040 996.000 371.320 1000.000 ;
    END
  END m_in[96]
  PIN m_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.180 996.000 375.460 1000.000 ;
    END
  END m_in[97]
  PIN m_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.860 996.000 379.140 1000.000 ;
    END
  END m_in[98]
  PIN m_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.540 996.000 382.820 1000.000 ;
    END
  END m_in[99]
  PIN m_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.240 996.000 35.520 1000.000 ;
    END
  END m_in[9]
  PIN m_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 3.440 998.810 4.040 ;
    END
  END m_out[0]
  PIN m_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 772.520 998.810 773.120 ;
    END
  END m_out[100]
  PIN m_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 780.000 998.810 780.600 ;
    END
  END m_out[101]
  PIN m_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 788.160 998.810 788.760 ;
    END
  END m_out[102]
  PIN m_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 795.640 998.810 796.240 ;
    END
  END m_out[103]
  PIN m_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 803.120 998.810 803.720 ;
    END
  END m_out[104]
  PIN m_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 811.280 998.810 811.880 ;
    END
  END m_out[105]
  PIN m_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 818.760 998.810 819.360 ;
    END
  END m_out[106]
  PIN m_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 826.240 998.810 826.840 ;
    END
  END m_out[107]
  PIN m_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 834.400 998.810 835.000 ;
    END
  END m_out[108]
  PIN m_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 841.880 998.810 842.480 ;
    END
  END m_out[109]
  PIN m_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 80.280 998.810 80.880 ;
    END
  END m_out[10]
  PIN m_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 849.360 998.810 849.960 ;
    END
  END m_out[110]
  PIN m_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 857.520 998.810 858.120 ;
    END
  END m_out[111]
  PIN m_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 865.000 998.810 865.600 ;
    END
  END m_out[112]
  PIN m_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 872.480 998.810 873.080 ;
    END
  END m_out[113]
  PIN m_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 879.960 998.810 880.560 ;
    END
  END m_out[114]
  PIN m_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 888.120 998.810 888.720 ;
    END
  END m_out[115]
  PIN m_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 895.600 998.810 896.200 ;
    END
  END m_out[116]
  PIN m_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 903.080 998.810 903.680 ;
    END
  END m_out[117]
  PIN m_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 911.240 998.810 911.840 ;
    END
  END m_out[118]
  PIN m_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 918.720 998.810 919.320 ;
    END
  END m_out[119]
  PIN m_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 87.760 998.810 88.360 ;
    END
  END m_out[11]
  PIN m_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 926.200 998.810 926.800 ;
    END
  END m_out[120]
  PIN m_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 934.360 998.810 934.960 ;
    END
  END m_out[121]
  PIN m_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 941.840 998.810 942.440 ;
    END
  END m_out[122]
  PIN m_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 949.320 998.810 949.920 ;
    END
  END m_out[123]
  PIN m_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 957.480 998.810 958.080 ;
    END
  END m_out[124]
  PIN m_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 964.960 998.810 965.560 ;
    END
  END m_out[125]
  PIN m_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 972.440 998.810 973.040 ;
    END
  END m_out[126]
  PIN m_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 980.600 998.810 981.200 ;
    END
  END m_out[127]
  PIN m_out[128]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 988.080 998.810 988.680 ;
    END
  END m_out[128]
  PIN m_out[129]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 995.560 998.810 996.160 ;
    END
  END m_out[129]
  PIN m_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 95.240 998.810 95.840 ;
    END
  END m_out[12]
  PIN m_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 103.400 998.810 104.000 ;
    END
  END m_out[13]
  PIN m_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 110.880 998.810 111.480 ;
    END
  END m_out[14]
  PIN m_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 118.360 998.810 118.960 ;
    END
  END m_out[15]
  PIN m_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 126.520 998.810 127.120 ;
    END
  END m_out[16]
  PIN m_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 134.000 998.810 134.600 ;
    END
  END m_out[17]
  PIN m_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 141.480 998.810 142.080 ;
    END
  END m_out[18]
  PIN m_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 148.960 998.810 149.560 ;
    END
  END m_out[19]
  PIN m_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 10.920 998.810 11.520 ;
    END
  END m_out[1]
  PIN m_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 157.120 998.810 157.720 ;
    END
  END m_out[20]
  PIN m_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 164.600 998.810 165.200 ;
    END
  END m_out[21]
  PIN m_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 172.080 998.810 172.680 ;
    END
  END m_out[22]
  PIN m_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 180.240 998.810 180.840 ;
    END
  END m_out[23]
  PIN m_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 187.720 998.810 188.320 ;
    END
  END m_out[24]
  PIN m_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 195.200 998.810 195.800 ;
    END
  END m_out[25]
  PIN m_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 203.360 998.810 203.960 ;
    END
  END m_out[26]
  PIN m_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 210.840 998.810 211.440 ;
    END
  END m_out[27]
  PIN m_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 218.320 998.810 218.920 ;
    END
  END m_out[28]
  PIN m_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 226.480 998.810 227.080 ;
    END
  END m_out[29]
  PIN m_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 18.400 998.810 19.000 ;
    END
  END m_out[2]
  PIN m_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 233.960 998.810 234.560 ;
    END
  END m_out[30]
  PIN m_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 241.440 998.810 242.040 ;
    END
  END m_out[31]
  PIN m_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 249.600 998.810 250.200 ;
    END
  END m_out[32]
  PIN m_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 257.080 998.810 257.680 ;
    END
  END m_out[33]
  PIN m_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 264.560 998.810 265.160 ;
    END
  END m_out[34]
  PIN m_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 272.720 998.810 273.320 ;
    END
  END m_out[35]
  PIN m_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 280.200 998.810 280.800 ;
    END
  END m_out[36]
  PIN m_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 287.680 998.810 288.280 ;
    END
  END m_out[37]
  PIN m_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 295.160 998.810 295.760 ;
    END
  END m_out[38]
  PIN m_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 303.320 998.810 303.920 ;
    END
  END m_out[39]
  PIN m_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 25.880 998.810 26.480 ;
    END
  END m_out[3]
  PIN m_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 310.800 998.810 311.400 ;
    END
  END m_out[40]
  PIN m_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 318.280 998.810 318.880 ;
    END
  END m_out[41]
  PIN m_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 326.440 998.810 327.040 ;
    END
  END m_out[42]
  PIN m_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 333.920 998.810 334.520 ;
    END
  END m_out[43]
  PIN m_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 341.400 998.810 342.000 ;
    END
  END m_out[44]
  PIN m_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 349.560 998.810 350.160 ;
    END
  END m_out[45]
  PIN m_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 357.040 998.810 357.640 ;
    END
  END m_out[46]
  PIN m_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 364.520 998.810 365.120 ;
    END
  END m_out[47]
  PIN m_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 372.680 998.810 373.280 ;
    END
  END m_out[48]
  PIN m_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 380.160 998.810 380.760 ;
    END
  END m_out[49]
  PIN m_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 34.040 998.810 34.640 ;
    END
  END m_out[4]
  PIN m_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 387.640 998.810 388.240 ;
    END
  END m_out[50]
  PIN m_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 395.800 998.810 396.400 ;
    END
  END m_out[51]
  PIN m_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 403.280 998.810 403.880 ;
    END
  END m_out[52]
  PIN m_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 410.760 998.810 411.360 ;
    END
  END m_out[53]
  PIN m_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 418.920 998.810 419.520 ;
    END
  END m_out[54]
  PIN m_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 426.400 998.810 427.000 ;
    END
  END m_out[55]
  PIN m_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 433.880 998.810 434.480 ;
    END
  END m_out[56]
  PIN m_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 441.360 998.810 441.960 ;
    END
  END m_out[57]
  PIN m_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 449.520 998.810 450.120 ;
    END
  END m_out[58]
  PIN m_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 457.000 998.810 457.600 ;
    END
  END m_out[59]
  PIN m_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 41.520 998.810 42.120 ;
    END
  END m_out[5]
  PIN m_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 464.480 998.810 465.080 ;
    END
  END m_out[60]
  PIN m_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 472.640 998.810 473.240 ;
    END
  END m_out[61]
  PIN m_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 480.120 998.810 480.720 ;
    END
  END m_out[62]
  PIN m_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 487.600 998.810 488.200 ;
    END
  END m_out[63]
  PIN m_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 495.760 998.810 496.360 ;
    END
  END m_out[64]
  PIN m_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 503.240 998.810 503.840 ;
    END
  END m_out[65]
  PIN m_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 510.720 998.810 511.320 ;
    END
  END m_out[66]
  PIN m_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 518.880 998.810 519.480 ;
    END
  END m_out[67]
  PIN m_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 526.360 998.810 526.960 ;
    END
  END m_out[68]
  PIN m_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 533.840 998.810 534.440 ;
    END
  END m_out[69]
  PIN m_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 49.000 998.810 49.600 ;
    END
  END m_out[6]
  PIN m_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 542.000 998.810 542.600 ;
    END
  END m_out[70]
  PIN m_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 549.480 998.810 550.080 ;
    END
  END m_out[71]
  PIN m_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 556.960 998.810 557.560 ;
    END
  END m_out[72]
  PIN m_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 565.120 998.810 565.720 ;
    END
  END m_out[73]
  PIN m_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 572.600 998.810 573.200 ;
    END
  END m_out[74]
  PIN m_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 580.080 998.810 580.680 ;
    END
  END m_out[75]
  PIN m_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 587.560 998.810 588.160 ;
    END
  END m_out[76]
  PIN m_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 595.720 998.810 596.320 ;
    END
  END m_out[77]
  PIN m_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 603.200 998.810 603.800 ;
    END
  END m_out[78]
  PIN m_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 610.680 998.810 611.280 ;
    END
  END m_out[79]
  PIN m_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 57.160 998.810 57.760 ;
    END
  END m_out[7]
  PIN m_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 618.840 998.810 619.440 ;
    END
  END m_out[80]
  PIN m_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 626.320 998.810 626.920 ;
    END
  END m_out[81]
  PIN m_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 633.800 998.810 634.400 ;
    END
  END m_out[82]
  PIN m_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 641.960 998.810 642.560 ;
    END
  END m_out[83]
  PIN m_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 649.440 998.810 650.040 ;
    END
  END m_out[84]
  PIN m_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 656.920 998.810 657.520 ;
    END
  END m_out[85]
  PIN m_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 665.080 998.810 665.680 ;
    END
  END m_out[86]
  PIN m_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 672.560 998.810 673.160 ;
    END
  END m_out[87]
  PIN m_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 680.040 998.810 680.640 ;
    END
  END m_out[88]
  PIN m_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 688.200 998.810 688.800 ;
    END
  END m_out[89]
  PIN m_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 64.640 998.810 65.240 ;
    END
  END m_out[8]
  PIN m_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 695.680 998.810 696.280 ;
    END
  END m_out[90]
  PIN m_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 703.160 998.810 703.760 ;
    END
  END m_out[91]
  PIN m_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 711.320 998.810 711.920 ;
    END
  END m_out[92]
  PIN m_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 718.800 998.810 719.400 ;
    END
  END m_out[93]
  PIN m_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 726.280 998.810 726.880 ;
    END
  END m_out[94]
  PIN m_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 733.760 998.810 734.360 ;
    END
  END m_out[95]
  PIN m_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 741.920 998.810 742.520 ;
    END
  END m_out[96]
  PIN m_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 749.400 998.810 750.000 ;
    END
  END m_out[97]
  PIN m_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 756.880 998.810 757.480 ;
    END
  END m_out[98]
  PIN m_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 765.040 998.810 765.640 ;
    END
  END m_out[99]
  PIN m_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 994.810 72.120 998.810 72.720 ;
    END
  END m_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 941.450 10.640 943.050 987.600 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 787.850 10.640 789.450 987.600 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 634.250 10.640 635.850 987.600 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 480.650 10.640 482.250 987.600 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 327.050 10.640 328.650 987.600 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 173.450 10.640 175.050 987.600 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.850 10.640 21.450 987.600 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 864.650 10.640 866.250 987.600 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 711.050 10.640 712.650 987.600 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 557.450 10.640 559.050 987.600 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 403.850 10.640 405.450 987.600 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 250.250 10.640 251.850 987.600 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.650 10.640 98.250 987.600 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 944.750 10.880 946.350 987.360 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 791.150 10.880 792.750 987.360 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 637.550 10.880 639.150 987.360 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 483.950 10.880 485.550 987.360 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 330.350 10.880 331.950 987.360 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 176.750 10.880 178.350 987.360 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 23.150 10.880 24.750 987.360 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 867.950 10.880 869.550 987.360 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 714.350 10.880 715.950 987.360 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 560.750 10.880 562.350 987.360 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 407.150 10.880 408.750 987.360 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 253.550 10.880 255.150 987.360 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 99.950 10.880 101.550 987.360 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 948.050 10.880 949.650 987.360 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 794.450 10.880 796.050 987.360 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 640.850 10.880 642.450 987.360 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 487.250 10.880 488.850 987.360 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 333.650 10.880 335.250 987.360 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 180.050 10.880 181.650 987.360 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 26.450 10.880 28.050 987.360 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 871.250 10.880 872.850 987.360 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 717.650 10.880 719.250 987.360 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 564.050 10.880 565.650 987.360 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 410.450 10.880 412.050 987.360 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 256.850 10.880 258.450 987.360 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 103.250 10.880 104.850 987.360 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 951.350 10.880 952.950 987.360 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 797.750 10.880 799.350 987.360 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 644.150 10.880 645.750 987.360 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 490.550 10.880 492.150 987.360 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 336.950 10.880 338.550 987.360 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 183.350 10.880 184.950 987.360 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 29.750 10.880 31.350 987.360 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 874.550 10.880 876.150 987.360 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 720.950 10.880 722.550 987.360 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 567.350 10.880 568.950 987.360 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 413.750 10.880 415.350 987.360 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 260.150 10.880 261.750 987.360 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 106.550 10.880 108.150 987.360 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 4.330 10.795 994.105 989.655 ;
      LAYER met1 ;
        RECT 0.720 1.740 996.940 999.900 ;
      LAYER met2 ;
        RECT 0.280 995.720 0.460 1000.125 ;
        RECT 1.300 995.720 4.140 1000.125 ;
        RECT 4.980 995.720 7.820 1000.125 ;
        RECT 8.660 995.720 11.960 1000.125 ;
        RECT 12.800 995.720 15.640 1000.125 ;
        RECT 16.480 995.720 19.320 1000.125 ;
        RECT 20.160 995.720 23.460 1000.125 ;
        RECT 24.300 995.720 27.140 1000.125 ;
        RECT 27.980 995.720 31.280 1000.125 ;
        RECT 32.120 995.720 34.960 1000.125 ;
        RECT 35.800 995.720 38.640 1000.125 ;
        RECT 39.480 995.720 42.780 1000.125 ;
        RECT 43.620 995.720 46.460 1000.125 ;
        RECT 47.300 995.720 50.600 1000.125 ;
        RECT 51.440 995.720 54.280 1000.125 ;
        RECT 55.120 995.720 57.960 1000.125 ;
        RECT 58.800 995.720 62.100 1000.125 ;
        RECT 62.940 995.720 65.780 1000.125 ;
        RECT 66.620 995.720 69.920 1000.125 ;
        RECT 70.760 995.720 73.600 1000.125 ;
        RECT 74.440 995.720 77.280 1000.125 ;
        RECT 78.120 995.720 81.420 1000.125 ;
        RECT 82.260 995.720 85.100 1000.125 ;
        RECT 85.940 995.720 89.240 1000.125 ;
        RECT 90.080 995.720 92.920 1000.125 ;
        RECT 93.760 995.720 96.600 1000.125 ;
        RECT 97.440 995.720 100.740 1000.125 ;
        RECT 101.580 995.720 104.420 1000.125 ;
        RECT 105.260 995.720 108.560 1000.125 ;
        RECT 109.400 995.720 112.240 1000.125 ;
        RECT 113.080 995.720 115.920 1000.125 ;
        RECT 116.760 995.720 120.060 1000.125 ;
        RECT 120.900 995.720 123.740 1000.125 ;
        RECT 124.580 995.720 127.420 1000.125 ;
        RECT 128.260 995.720 131.560 1000.125 ;
        RECT 132.400 995.720 135.240 1000.125 ;
        RECT 136.080 995.720 139.380 1000.125 ;
        RECT 140.220 995.720 143.060 1000.125 ;
        RECT 143.900 995.720 146.740 1000.125 ;
        RECT 147.580 995.720 150.880 1000.125 ;
        RECT 151.720 995.720 154.560 1000.125 ;
        RECT 155.400 995.720 158.700 1000.125 ;
        RECT 159.540 995.720 162.380 1000.125 ;
        RECT 163.220 995.720 166.060 1000.125 ;
        RECT 166.900 995.720 170.200 1000.125 ;
        RECT 171.040 995.720 173.880 1000.125 ;
        RECT 174.720 995.720 178.020 1000.125 ;
        RECT 178.860 995.720 181.700 1000.125 ;
        RECT 182.540 995.720 185.380 1000.125 ;
        RECT 186.220 995.720 189.520 1000.125 ;
        RECT 190.360 995.720 193.200 1000.125 ;
        RECT 194.040 995.720 197.340 1000.125 ;
        RECT 198.180 995.720 201.020 1000.125 ;
        RECT 201.860 995.720 204.700 1000.125 ;
        RECT 205.540 995.720 208.840 1000.125 ;
        RECT 209.680 995.720 212.520 1000.125 ;
        RECT 213.360 995.720 216.660 1000.125 ;
        RECT 217.500 995.720 220.340 1000.125 ;
        RECT 221.180 995.720 224.020 1000.125 ;
        RECT 224.860 995.720 228.160 1000.125 ;
        RECT 229.000 995.720 231.840 1000.125 ;
        RECT 232.680 995.720 235.980 1000.125 ;
        RECT 236.820 995.720 239.660 1000.125 ;
        RECT 240.500 995.720 243.340 1000.125 ;
        RECT 244.180 995.720 247.480 1000.125 ;
        RECT 248.320 995.720 251.160 1000.125 ;
        RECT 252.000 995.720 254.840 1000.125 ;
        RECT 255.680 995.720 258.980 1000.125 ;
        RECT 259.820 995.720 262.660 1000.125 ;
        RECT 263.500 995.720 266.800 1000.125 ;
        RECT 267.640 995.720 270.480 1000.125 ;
        RECT 271.320 995.720 274.160 1000.125 ;
        RECT 275.000 995.720 278.300 1000.125 ;
        RECT 279.140 995.720 281.980 1000.125 ;
        RECT 282.820 995.720 286.120 1000.125 ;
        RECT 286.960 995.720 289.800 1000.125 ;
        RECT 290.640 995.720 293.480 1000.125 ;
        RECT 294.320 995.720 297.620 1000.125 ;
        RECT 298.460 995.720 301.300 1000.125 ;
        RECT 302.140 995.720 305.440 1000.125 ;
        RECT 306.280 995.720 309.120 1000.125 ;
        RECT 309.960 995.720 312.800 1000.125 ;
        RECT 313.640 995.720 316.940 1000.125 ;
        RECT 317.780 995.720 320.620 1000.125 ;
        RECT 321.460 995.720 324.760 1000.125 ;
        RECT 325.600 995.720 328.440 1000.125 ;
        RECT 329.280 995.720 332.120 1000.125 ;
        RECT 332.960 995.720 336.260 1000.125 ;
        RECT 337.100 995.720 339.940 1000.125 ;
        RECT 340.780 995.720 344.080 1000.125 ;
        RECT 344.920 995.720 347.760 1000.125 ;
        RECT 348.600 995.720 351.440 1000.125 ;
        RECT 352.280 995.720 355.580 1000.125 ;
        RECT 356.420 995.720 359.260 1000.125 ;
        RECT 360.100 995.720 363.400 1000.125 ;
        RECT 364.240 995.720 367.080 1000.125 ;
        RECT 367.920 995.720 370.760 1000.125 ;
        RECT 371.600 995.720 374.900 1000.125 ;
        RECT 375.740 995.720 378.580 1000.125 ;
        RECT 379.420 995.720 382.260 1000.125 ;
        RECT 383.100 995.720 386.400 1000.125 ;
        RECT 387.240 995.720 390.080 1000.125 ;
        RECT 390.920 995.720 394.220 1000.125 ;
        RECT 395.060 995.720 397.900 1000.125 ;
        RECT 398.740 995.720 401.580 1000.125 ;
        RECT 402.420 995.720 405.720 1000.125 ;
        RECT 406.560 995.720 409.400 1000.125 ;
        RECT 410.240 995.720 413.540 1000.125 ;
        RECT 414.380 995.720 417.220 1000.125 ;
        RECT 418.060 995.720 420.900 1000.125 ;
        RECT 421.740 995.720 425.040 1000.125 ;
        RECT 425.880 995.720 428.720 1000.125 ;
        RECT 429.560 995.720 432.860 1000.125 ;
        RECT 433.700 995.720 436.540 1000.125 ;
        RECT 437.380 995.720 440.220 1000.125 ;
        RECT 441.060 995.720 444.360 1000.125 ;
        RECT 445.200 995.720 448.040 1000.125 ;
        RECT 448.880 995.720 452.180 1000.125 ;
        RECT 453.020 995.720 455.860 1000.125 ;
        RECT 456.700 995.720 459.540 1000.125 ;
        RECT 460.380 995.720 463.680 1000.125 ;
        RECT 464.520 995.720 467.360 1000.125 ;
        RECT 468.200 995.720 471.500 1000.125 ;
        RECT 472.340 995.720 475.180 1000.125 ;
        RECT 476.020 995.720 478.860 1000.125 ;
        RECT 479.700 995.720 483.000 1000.125 ;
        RECT 483.840 995.720 486.680 1000.125 ;
        RECT 487.520 995.720 490.820 1000.125 ;
        RECT 491.660 995.720 494.500 1000.125 ;
        RECT 495.340 995.720 498.180 1000.125 ;
        RECT 499.020 995.720 502.320 1000.125 ;
        RECT 503.160 995.720 506.000 1000.125 ;
        RECT 506.840 995.720 509.680 1000.125 ;
        RECT 510.520 995.720 513.820 1000.125 ;
        RECT 514.660 995.720 517.500 1000.125 ;
        RECT 518.340 995.720 521.640 1000.125 ;
        RECT 522.480 995.720 525.320 1000.125 ;
        RECT 526.160 995.720 529.000 1000.125 ;
        RECT 529.840 995.720 533.140 1000.125 ;
        RECT 533.980 995.720 536.820 1000.125 ;
        RECT 537.660 995.720 540.960 1000.125 ;
        RECT 541.800 995.720 544.640 1000.125 ;
        RECT 545.480 995.720 548.320 1000.125 ;
        RECT 549.160 995.720 552.460 1000.125 ;
        RECT 553.300 995.720 556.140 1000.125 ;
        RECT 556.980 995.720 560.280 1000.125 ;
        RECT 561.120 995.720 563.960 1000.125 ;
        RECT 564.800 995.720 567.640 1000.125 ;
        RECT 568.480 995.720 571.780 1000.125 ;
        RECT 572.620 995.720 575.460 1000.125 ;
        RECT 576.300 995.720 579.600 1000.125 ;
        RECT 580.440 995.720 583.280 1000.125 ;
        RECT 584.120 995.720 586.960 1000.125 ;
        RECT 587.800 995.720 591.100 1000.125 ;
        RECT 591.940 995.720 594.780 1000.125 ;
        RECT 595.620 995.720 598.920 1000.125 ;
        RECT 599.760 995.720 602.600 1000.125 ;
        RECT 603.440 995.720 606.280 1000.125 ;
        RECT 607.120 995.720 610.420 1000.125 ;
        RECT 611.260 995.720 614.100 1000.125 ;
        RECT 614.940 995.720 618.240 1000.125 ;
        RECT 619.080 995.720 621.920 1000.125 ;
        RECT 622.760 995.720 625.600 1000.125 ;
        RECT 626.440 995.720 629.740 1000.125 ;
        RECT 630.580 995.720 633.420 1000.125 ;
        RECT 634.260 995.720 637.100 1000.125 ;
        RECT 637.940 995.720 641.240 1000.125 ;
        RECT 642.080 995.720 644.920 1000.125 ;
        RECT 645.760 995.720 649.060 1000.125 ;
        RECT 649.900 995.720 652.740 1000.125 ;
        RECT 653.580 995.720 656.420 1000.125 ;
        RECT 657.260 995.720 660.560 1000.125 ;
        RECT 661.400 995.720 664.240 1000.125 ;
        RECT 665.080 995.720 668.380 1000.125 ;
        RECT 669.220 995.720 672.060 1000.125 ;
        RECT 672.900 995.720 675.740 1000.125 ;
        RECT 676.580 995.720 679.880 1000.125 ;
        RECT 680.720 995.720 683.560 1000.125 ;
        RECT 684.400 995.720 687.700 1000.125 ;
        RECT 688.540 995.720 691.380 1000.125 ;
        RECT 692.220 995.720 695.060 1000.125 ;
        RECT 695.900 995.720 699.200 1000.125 ;
        RECT 700.040 995.720 702.880 1000.125 ;
        RECT 703.720 995.720 707.020 1000.125 ;
        RECT 707.860 995.720 710.700 1000.125 ;
        RECT 711.540 995.720 714.380 1000.125 ;
        RECT 715.220 995.720 718.520 1000.125 ;
        RECT 719.360 995.720 722.200 1000.125 ;
        RECT 723.040 995.720 726.340 1000.125 ;
        RECT 727.180 995.720 730.020 1000.125 ;
        RECT 730.860 995.720 733.700 1000.125 ;
        RECT 734.540 995.720 737.840 1000.125 ;
        RECT 738.680 995.720 741.520 1000.125 ;
        RECT 742.360 995.720 745.660 1000.125 ;
        RECT 746.500 995.720 749.340 1000.125 ;
        RECT 750.180 995.720 753.020 1000.125 ;
        RECT 753.860 995.720 757.160 1000.125 ;
        RECT 758.000 995.720 760.840 1000.125 ;
        RECT 761.680 995.720 764.520 1000.125 ;
        RECT 765.360 995.720 768.660 1000.125 ;
        RECT 769.500 995.720 772.340 1000.125 ;
        RECT 773.180 995.720 776.480 1000.125 ;
        RECT 777.320 995.720 780.160 1000.125 ;
        RECT 781.000 995.720 783.840 1000.125 ;
        RECT 784.680 995.720 787.980 1000.125 ;
        RECT 788.820 995.720 791.660 1000.125 ;
        RECT 792.500 995.720 795.800 1000.125 ;
        RECT 796.640 995.720 799.480 1000.125 ;
        RECT 800.320 995.720 803.160 1000.125 ;
        RECT 804.000 995.720 807.300 1000.125 ;
        RECT 808.140 995.720 810.980 1000.125 ;
        RECT 811.820 995.720 815.120 1000.125 ;
        RECT 815.960 995.720 818.800 1000.125 ;
        RECT 819.640 995.720 822.480 1000.125 ;
        RECT 823.320 995.720 826.620 1000.125 ;
        RECT 827.460 995.720 830.300 1000.125 ;
        RECT 831.140 995.720 834.440 1000.125 ;
        RECT 835.280 995.720 838.120 1000.125 ;
        RECT 838.960 995.720 841.800 1000.125 ;
        RECT 842.640 995.720 845.940 1000.125 ;
        RECT 846.780 995.720 849.620 1000.125 ;
        RECT 850.460 995.720 853.760 1000.125 ;
        RECT 854.600 995.720 857.440 1000.125 ;
        RECT 858.280 995.720 861.120 1000.125 ;
        RECT 861.960 995.720 865.260 1000.125 ;
        RECT 866.100 995.720 868.940 1000.125 ;
        RECT 869.780 995.720 873.080 1000.125 ;
        RECT 873.920 995.720 876.760 1000.125 ;
        RECT 877.600 995.720 880.440 1000.125 ;
        RECT 881.280 995.720 884.580 1000.125 ;
        RECT 885.420 995.720 888.260 1000.125 ;
        RECT 889.100 995.720 891.940 1000.125 ;
        RECT 892.780 995.720 896.080 1000.125 ;
        RECT 896.920 995.720 899.760 1000.125 ;
        RECT 900.600 995.720 903.900 1000.125 ;
        RECT 904.740 995.720 907.580 1000.125 ;
        RECT 908.420 995.720 911.260 1000.125 ;
        RECT 912.100 995.720 915.400 1000.125 ;
        RECT 916.240 995.720 919.080 1000.125 ;
        RECT 919.920 995.720 923.220 1000.125 ;
        RECT 924.060 995.720 926.900 1000.125 ;
        RECT 927.740 995.720 930.580 1000.125 ;
        RECT 931.420 995.720 934.720 1000.125 ;
        RECT 935.560 995.720 938.400 1000.125 ;
        RECT 939.240 995.720 942.540 1000.125 ;
        RECT 943.380 995.720 946.220 1000.125 ;
        RECT 947.060 995.720 949.900 1000.125 ;
        RECT 950.740 995.720 954.040 1000.125 ;
        RECT 954.880 995.720 957.720 1000.125 ;
        RECT 958.560 995.720 961.860 1000.125 ;
        RECT 962.700 995.720 965.540 1000.125 ;
        RECT 966.380 995.720 969.220 1000.125 ;
        RECT 970.060 995.720 973.360 1000.125 ;
        RECT 974.200 995.720 977.040 1000.125 ;
        RECT 977.880 995.720 981.180 1000.125 ;
        RECT 982.020 995.720 984.860 1000.125 ;
        RECT 985.700 995.720 988.540 1000.125 ;
        RECT 989.380 995.720 992.680 1000.125 ;
        RECT 993.520 995.720 996.360 1000.125 ;
        RECT 0.280 4.280 996.910 995.720 ;
        RECT 0.280 1.710 498.640 4.280 ;
        RECT 499.480 1.710 996.910 4.280 ;
      LAYER met3 ;
        RECT 0.000 996.560 995.105 1000.105 ;
        RECT 0.000 995.160 994.410 996.560 ;
        RECT 0.000 989.080 995.105 995.160 ;
        RECT 0.000 987.680 994.410 989.080 ;
        RECT 0.000 981.600 995.105 987.680 ;
        RECT 0.000 980.200 994.410 981.600 ;
        RECT 0.000 973.440 995.105 980.200 ;
        RECT 0.000 972.040 994.410 973.440 ;
        RECT 0.000 965.960 995.105 972.040 ;
        RECT 0.000 964.560 994.410 965.960 ;
        RECT 0.000 958.480 995.105 964.560 ;
        RECT 0.000 957.080 994.410 958.480 ;
        RECT 0.000 950.320 995.105 957.080 ;
        RECT 0.000 948.920 994.410 950.320 ;
        RECT 0.000 942.840 995.105 948.920 ;
        RECT 0.000 941.440 994.410 942.840 ;
        RECT 0.000 935.360 995.105 941.440 ;
        RECT 0.000 933.960 994.410 935.360 ;
        RECT 0.000 927.200 995.105 933.960 ;
        RECT 0.000 925.800 994.410 927.200 ;
        RECT 0.000 919.720 995.105 925.800 ;
        RECT 0.000 918.320 994.410 919.720 ;
        RECT 0.000 912.240 995.105 918.320 ;
        RECT 0.000 910.840 994.410 912.240 ;
        RECT 0.000 904.080 995.105 910.840 ;
        RECT 0.000 902.680 994.410 904.080 ;
        RECT 0.000 896.600 995.105 902.680 ;
        RECT 0.000 895.200 994.410 896.600 ;
        RECT 0.000 889.120 995.105 895.200 ;
        RECT 0.000 887.720 994.410 889.120 ;
        RECT 0.000 880.960 995.105 887.720 ;
        RECT 0.000 879.560 994.410 880.960 ;
        RECT 0.000 873.480 995.105 879.560 ;
        RECT 0.000 872.080 994.410 873.480 ;
        RECT 0.000 866.000 995.105 872.080 ;
        RECT 0.000 864.600 994.410 866.000 ;
        RECT 0.000 858.520 995.105 864.600 ;
        RECT 0.000 857.120 994.410 858.520 ;
        RECT 0.000 850.360 995.105 857.120 ;
        RECT 0.000 848.960 994.410 850.360 ;
        RECT 0.000 842.880 995.105 848.960 ;
        RECT 0.000 841.480 994.410 842.880 ;
        RECT 0.000 835.400 995.105 841.480 ;
        RECT 0.000 834.000 994.410 835.400 ;
        RECT 0.000 827.240 995.105 834.000 ;
        RECT 0.000 825.840 994.410 827.240 ;
        RECT 0.000 819.760 995.105 825.840 ;
        RECT 0.000 818.360 994.410 819.760 ;
        RECT 0.000 812.280 995.105 818.360 ;
        RECT 0.000 810.880 994.410 812.280 ;
        RECT 0.000 804.120 995.105 810.880 ;
        RECT 0.000 802.720 994.410 804.120 ;
        RECT 0.000 796.640 995.105 802.720 ;
        RECT 0.000 795.240 994.410 796.640 ;
        RECT 0.000 789.160 995.105 795.240 ;
        RECT 0.000 787.760 994.410 789.160 ;
        RECT 0.000 781.000 995.105 787.760 ;
        RECT 0.000 779.600 994.410 781.000 ;
        RECT 0.000 773.520 995.105 779.600 ;
        RECT 0.000 772.120 994.410 773.520 ;
        RECT 0.000 766.040 995.105 772.120 ;
        RECT 0.000 764.640 994.410 766.040 ;
        RECT 0.000 757.880 995.105 764.640 ;
        RECT 0.000 756.480 994.410 757.880 ;
        RECT 0.000 750.400 995.105 756.480 ;
        RECT 0.000 749.000 994.410 750.400 ;
        RECT 0.000 742.920 995.105 749.000 ;
        RECT 0.000 741.520 994.410 742.920 ;
        RECT 0.000 734.760 995.105 741.520 ;
        RECT 0.000 733.360 994.410 734.760 ;
        RECT 0.000 727.280 995.105 733.360 ;
        RECT 0.000 725.880 994.410 727.280 ;
        RECT 0.000 719.800 995.105 725.880 ;
        RECT 0.000 718.400 994.410 719.800 ;
        RECT 0.000 712.320 995.105 718.400 ;
        RECT 0.000 710.920 994.410 712.320 ;
        RECT 0.000 704.160 995.105 710.920 ;
        RECT 0.000 702.760 994.410 704.160 ;
        RECT 0.000 696.680 995.105 702.760 ;
        RECT 0.000 695.280 994.410 696.680 ;
        RECT 0.000 689.200 995.105 695.280 ;
        RECT 0.000 687.800 994.410 689.200 ;
        RECT 0.000 681.040 995.105 687.800 ;
        RECT 0.000 679.640 994.410 681.040 ;
        RECT 0.000 673.560 995.105 679.640 ;
        RECT 0.000 672.160 994.410 673.560 ;
        RECT 0.000 666.080 995.105 672.160 ;
        RECT 0.000 664.680 994.410 666.080 ;
        RECT 0.000 657.920 995.105 664.680 ;
        RECT 0.000 656.520 994.410 657.920 ;
        RECT 0.000 650.440 995.105 656.520 ;
        RECT 0.000 649.040 994.410 650.440 ;
        RECT 0.000 642.960 995.105 649.040 ;
        RECT 0.000 641.560 994.410 642.960 ;
        RECT 0.000 634.800 995.105 641.560 ;
        RECT 0.000 633.400 994.410 634.800 ;
        RECT 0.000 627.320 995.105 633.400 ;
        RECT 0.000 625.920 994.410 627.320 ;
        RECT 0.000 619.840 995.105 625.920 ;
        RECT 0.000 618.440 994.410 619.840 ;
        RECT 0.000 611.680 995.105 618.440 ;
        RECT 0.000 610.280 994.410 611.680 ;
        RECT 0.000 604.200 995.105 610.280 ;
        RECT 0.000 602.800 994.410 604.200 ;
        RECT 0.000 596.720 995.105 602.800 ;
        RECT 0.000 595.320 994.410 596.720 ;
        RECT 0.000 588.560 995.105 595.320 ;
        RECT 0.000 587.160 994.410 588.560 ;
        RECT 0.000 581.080 995.105 587.160 ;
        RECT 0.000 579.680 994.410 581.080 ;
        RECT 0.000 573.600 995.105 579.680 ;
        RECT 0.000 572.200 994.410 573.600 ;
        RECT 0.000 566.120 995.105 572.200 ;
        RECT 0.000 564.720 994.410 566.120 ;
        RECT 0.000 557.960 995.105 564.720 ;
        RECT 0.000 556.560 994.410 557.960 ;
        RECT 0.000 550.480 995.105 556.560 ;
        RECT 0.000 549.080 994.410 550.480 ;
        RECT 0.000 543.000 995.105 549.080 ;
        RECT 0.000 541.600 994.410 543.000 ;
        RECT 0.000 534.840 995.105 541.600 ;
        RECT 0.000 533.440 994.410 534.840 ;
        RECT 0.000 527.360 995.105 533.440 ;
        RECT 0.000 525.960 994.410 527.360 ;
        RECT 0.000 519.880 995.105 525.960 ;
        RECT 0.000 518.480 994.410 519.880 ;
        RECT 0.000 511.720 995.105 518.480 ;
        RECT 0.000 510.320 994.410 511.720 ;
        RECT 0.000 504.240 995.105 510.320 ;
        RECT 0.000 502.840 994.410 504.240 ;
        RECT 0.000 496.760 995.105 502.840 ;
        RECT 0.000 495.360 994.410 496.760 ;
        RECT 0.000 488.600 995.105 495.360 ;
        RECT 0.000 487.200 994.410 488.600 ;
        RECT 0.000 481.120 995.105 487.200 ;
        RECT 0.000 479.720 994.410 481.120 ;
        RECT 0.000 473.640 995.105 479.720 ;
        RECT 0.000 472.240 994.410 473.640 ;
        RECT 0.000 465.480 995.105 472.240 ;
        RECT 0.000 464.080 994.410 465.480 ;
        RECT 0.000 458.000 995.105 464.080 ;
        RECT 0.000 456.600 994.410 458.000 ;
        RECT 0.000 450.520 995.105 456.600 ;
        RECT 0.000 449.120 994.410 450.520 ;
        RECT 0.000 442.360 995.105 449.120 ;
        RECT 0.000 440.960 994.410 442.360 ;
        RECT 0.000 434.880 995.105 440.960 ;
        RECT 0.000 433.480 994.410 434.880 ;
        RECT 0.000 427.400 995.105 433.480 ;
        RECT 0.000 426.000 994.410 427.400 ;
        RECT 0.000 419.920 995.105 426.000 ;
        RECT 0.000 418.520 994.410 419.920 ;
        RECT 0.000 411.760 995.105 418.520 ;
        RECT 0.000 410.360 994.410 411.760 ;
        RECT 0.000 404.280 995.105 410.360 ;
        RECT 0.000 402.880 994.410 404.280 ;
        RECT 0.000 396.800 995.105 402.880 ;
        RECT 0.000 395.400 994.410 396.800 ;
        RECT 0.000 388.640 995.105 395.400 ;
        RECT 0.000 387.240 994.410 388.640 ;
        RECT 0.000 381.160 995.105 387.240 ;
        RECT 0.000 379.760 994.410 381.160 ;
        RECT 0.000 373.680 995.105 379.760 ;
        RECT 0.000 372.280 994.410 373.680 ;
        RECT 0.000 365.520 995.105 372.280 ;
        RECT 0.000 364.120 994.410 365.520 ;
        RECT 0.000 358.040 995.105 364.120 ;
        RECT 0.000 356.640 994.410 358.040 ;
        RECT 0.000 350.560 995.105 356.640 ;
        RECT 0.000 349.160 994.410 350.560 ;
        RECT 0.000 342.400 995.105 349.160 ;
        RECT 0.000 341.000 994.410 342.400 ;
        RECT 0.000 334.920 995.105 341.000 ;
        RECT 0.000 333.520 994.410 334.920 ;
        RECT 0.000 327.440 995.105 333.520 ;
        RECT 0.000 326.040 994.410 327.440 ;
        RECT 0.000 319.280 995.105 326.040 ;
        RECT 0.000 317.880 994.410 319.280 ;
        RECT 0.000 311.800 995.105 317.880 ;
        RECT 0.000 310.400 994.410 311.800 ;
        RECT 0.000 304.320 995.105 310.400 ;
        RECT 0.000 302.920 994.410 304.320 ;
        RECT 0.000 296.160 995.105 302.920 ;
        RECT 0.000 294.760 994.410 296.160 ;
        RECT 0.000 288.680 995.105 294.760 ;
        RECT 0.000 287.280 994.410 288.680 ;
        RECT 0.000 281.200 995.105 287.280 ;
        RECT 0.000 279.800 994.410 281.200 ;
        RECT 0.000 273.720 995.105 279.800 ;
        RECT 0.000 272.320 994.410 273.720 ;
        RECT 0.000 265.560 995.105 272.320 ;
        RECT 0.000 264.160 994.410 265.560 ;
        RECT 0.000 258.080 995.105 264.160 ;
        RECT 0.000 256.680 994.410 258.080 ;
        RECT 0.000 250.600 995.105 256.680 ;
        RECT 0.000 249.200 994.410 250.600 ;
        RECT 0.000 242.440 995.105 249.200 ;
        RECT 0.000 241.040 994.410 242.440 ;
        RECT 0.000 234.960 995.105 241.040 ;
        RECT 0.000 233.560 994.410 234.960 ;
        RECT 0.000 227.480 995.105 233.560 ;
        RECT 0.000 226.080 994.410 227.480 ;
        RECT 0.000 219.320 995.105 226.080 ;
        RECT 0.000 217.920 994.410 219.320 ;
        RECT 0.000 211.840 995.105 217.920 ;
        RECT 0.000 210.440 994.410 211.840 ;
        RECT 0.000 204.360 995.105 210.440 ;
        RECT 0.000 202.960 994.410 204.360 ;
        RECT 0.000 196.200 995.105 202.960 ;
        RECT 0.000 194.800 994.410 196.200 ;
        RECT 0.000 188.720 995.105 194.800 ;
        RECT 0.000 187.320 994.410 188.720 ;
        RECT 0.000 181.240 995.105 187.320 ;
        RECT 0.000 179.840 994.410 181.240 ;
        RECT 0.000 173.080 995.105 179.840 ;
        RECT 0.000 171.680 994.410 173.080 ;
        RECT 0.000 165.600 995.105 171.680 ;
        RECT 0.000 164.200 994.410 165.600 ;
        RECT 0.000 158.120 995.105 164.200 ;
        RECT 0.000 156.720 994.410 158.120 ;
        RECT 0.000 149.960 995.105 156.720 ;
        RECT 0.000 148.560 994.410 149.960 ;
        RECT 0.000 142.480 995.105 148.560 ;
        RECT 0.000 141.080 994.410 142.480 ;
        RECT 0.000 135.000 995.105 141.080 ;
        RECT 0.000 133.600 994.410 135.000 ;
        RECT 0.000 127.520 995.105 133.600 ;
        RECT 0.000 126.120 994.410 127.520 ;
        RECT 0.000 119.360 995.105 126.120 ;
        RECT 0.000 117.960 994.410 119.360 ;
        RECT 0.000 111.880 995.105 117.960 ;
        RECT 0.000 110.480 994.410 111.880 ;
        RECT 0.000 104.400 995.105 110.480 ;
        RECT 0.000 103.000 994.410 104.400 ;
        RECT 0.000 96.240 995.105 103.000 ;
        RECT 0.000 94.840 994.410 96.240 ;
        RECT 0.000 88.760 995.105 94.840 ;
        RECT 0.000 87.360 994.410 88.760 ;
        RECT 0.000 81.280 995.105 87.360 ;
        RECT 0.000 79.880 994.410 81.280 ;
        RECT 0.000 73.120 995.105 79.880 ;
        RECT 0.000 71.720 994.410 73.120 ;
        RECT 0.000 65.640 995.105 71.720 ;
        RECT 0.000 64.240 994.410 65.640 ;
        RECT 0.000 58.160 995.105 64.240 ;
        RECT 0.000 56.760 994.410 58.160 ;
        RECT 0.000 50.000 995.105 56.760 ;
        RECT 0.000 48.600 994.410 50.000 ;
        RECT 0.000 42.520 995.105 48.600 ;
        RECT 0.000 41.120 994.410 42.520 ;
        RECT 0.000 35.040 995.105 41.120 ;
        RECT 0.000 33.640 994.410 35.040 ;
        RECT 0.000 26.880 995.105 33.640 ;
        RECT 0.000 25.480 994.410 26.880 ;
        RECT 0.000 19.400 995.105 25.480 ;
        RECT 0.000 18.000 994.410 19.400 ;
        RECT 0.000 11.920 995.105 18.000 ;
        RECT 0.000 10.520 994.410 11.920 ;
        RECT 0.000 4.440 995.105 10.520 ;
        RECT 0.000 3.040 994.410 4.440 ;
        RECT 0.000 2.895 995.105 3.040 ;
      LAYER met4 ;
        RECT 0.025 988.000 984.755 989.905 ;
        RECT 0.025 10.240 19.450 988.000 ;
        RECT 21.850 987.760 96.250 988.000 ;
        RECT 21.850 10.480 22.750 987.760 ;
        RECT 25.150 10.480 26.050 987.760 ;
        RECT 28.450 10.480 29.350 987.760 ;
        RECT 31.750 10.480 96.250 987.760 ;
        RECT 21.850 10.240 96.250 10.480 ;
        RECT 98.650 987.760 173.050 988.000 ;
        RECT 98.650 10.480 99.550 987.760 ;
        RECT 101.950 10.480 102.850 987.760 ;
        RECT 105.250 10.480 106.150 987.760 ;
        RECT 108.550 10.480 173.050 987.760 ;
        RECT 98.650 10.240 173.050 10.480 ;
        RECT 175.450 987.760 249.850 988.000 ;
        RECT 175.450 10.480 176.350 987.760 ;
        RECT 178.750 10.480 179.650 987.760 ;
        RECT 182.050 10.480 182.950 987.760 ;
        RECT 185.350 10.480 249.850 987.760 ;
        RECT 175.450 10.240 249.850 10.480 ;
        RECT 252.250 987.760 326.650 988.000 ;
        RECT 252.250 10.480 253.150 987.760 ;
        RECT 255.550 10.480 256.450 987.760 ;
        RECT 258.850 10.480 259.750 987.760 ;
        RECT 262.150 10.480 326.650 987.760 ;
        RECT 252.250 10.240 326.650 10.480 ;
        RECT 329.050 987.760 403.450 988.000 ;
        RECT 329.050 10.480 329.950 987.760 ;
        RECT 332.350 10.480 333.250 987.760 ;
        RECT 335.650 10.480 336.550 987.760 ;
        RECT 338.950 10.480 403.450 987.760 ;
        RECT 329.050 10.240 403.450 10.480 ;
        RECT 405.850 987.760 480.250 988.000 ;
        RECT 405.850 10.480 406.750 987.760 ;
        RECT 409.150 10.480 410.050 987.760 ;
        RECT 412.450 10.480 413.350 987.760 ;
        RECT 415.750 10.480 480.250 987.760 ;
        RECT 405.850 10.240 480.250 10.480 ;
        RECT 482.650 987.760 557.050 988.000 ;
        RECT 482.650 10.480 483.550 987.760 ;
        RECT 485.950 10.480 486.850 987.760 ;
        RECT 489.250 10.480 490.150 987.760 ;
        RECT 492.550 10.480 557.050 987.760 ;
        RECT 482.650 10.240 557.050 10.480 ;
        RECT 559.450 987.760 633.850 988.000 ;
        RECT 559.450 10.480 560.350 987.760 ;
        RECT 562.750 10.480 563.650 987.760 ;
        RECT 566.050 10.480 566.950 987.760 ;
        RECT 569.350 10.480 633.850 987.760 ;
        RECT 559.450 10.240 633.850 10.480 ;
        RECT 636.250 987.760 710.650 988.000 ;
        RECT 636.250 10.480 637.150 987.760 ;
        RECT 639.550 10.480 640.450 987.760 ;
        RECT 642.850 10.480 643.750 987.760 ;
        RECT 646.150 10.480 710.650 987.760 ;
        RECT 636.250 10.240 710.650 10.480 ;
        RECT 713.050 987.760 787.450 988.000 ;
        RECT 713.050 10.480 713.950 987.760 ;
        RECT 716.350 10.480 717.250 987.760 ;
        RECT 719.650 10.480 720.550 987.760 ;
        RECT 722.950 10.480 787.450 987.760 ;
        RECT 713.050 10.240 787.450 10.480 ;
        RECT 789.850 987.760 864.250 988.000 ;
        RECT 789.850 10.480 790.750 987.760 ;
        RECT 793.150 10.480 794.050 987.760 ;
        RECT 796.450 10.480 797.350 987.760 ;
        RECT 799.750 10.480 864.250 987.760 ;
        RECT 789.850 10.240 864.250 10.480 ;
        RECT 866.650 987.760 941.050 988.000 ;
        RECT 866.650 10.480 867.550 987.760 ;
        RECT 869.950 10.480 870.850 987.760 ;
        RECT 873.250 10.480 874.150 987.760 ;
        RECT 876.550 10.480 941.050 987.760 ;
        RECT 866.650 10.240 941.050 10.480 ;
        RECT 943.450 987.760 984.755 988.000 ;
        RECT 943.450 10.480 944.350 987.760 ;
        RECT 946.750 10.480 947.650 987.760 ;
        RECT 950.050 10.480 950.950 987.760 ;
        RECT 953.350 10.480 984.755 987.760 ;
        RECT 943.450 10.240 984.755 10.480 ;
        RECT 0.025 2.895 984.755 10.240 ;
  END
END multiply_4
END LIBRARY

