magic
tech sky130A
magscale 1 2
timestamp 1608844368
<< obsli1 >>
rect 814 1607 158749 158279
<< obsm1 >>
rect 0 1088 159408 158288
<< metal2 >>
rect 4 158648 60 159448
rect 556 158648 612 159448
rect 1200 158648 1256 159448
rect 1844 158648 1900 159448
rect 2396 158648 2452 159448
rect 3040 158648 3096 159448
rect 3684 158648 3740 159448
rect 4236 158648 4292 159448
rect 4880 158648 4936 159448
rect 5524 158648 5580 159448
rect 6076 158648 6132 159448
rect 6720 158648 6776 159448
rect 7364 158648 7420 159448
rect 7916 158648 7972 159448
rect 8560 158648 8616 159448
rect 9204 158648 9260 159448
rect 9848 158648 9904 159448
rect 10400 158648 10456 159448
rect 11044 158648 11100 159448
rect 11688 158648 11744 159448
rect 12240 158648 12296 159448
rect 12884 158648 12940 159448
rect 13528 158648 13584 159448
rect 14080 158648 14136 159448
rect 14724 158648 14780 159448
rect 15368 158648 15424 159448
rect 15920 158648 15976 159448
rect 16564 158648 16620 159448
rect 17208 158648 17264 159448
rect 17760 158648 17816 159448
rect 18404 158648 18460 159448
rect 19048 158648 19104 159448
rect 19692 158648 19748 159448
rect 20244 158648 20300 159448
rect 20888 158648 20944 159448
rect 21532 158648 21588 159448
rect 22084 158648 22140 159448
rect 22728 158648 22784 159448
rect 23372 158648 23428 159448
rect 23924 158648 23980 159448
rect 24568 158648 24624 159448
rect 25212 158648 25268 159448
rect 25764 158648 25820 159448
rect 26408 158648 26464 159448
rect 27052 158648 27108 159448
rect 27604 158648 27660 159448
rect 28248 158648 28304 159448
rect 28892 158648 28948 159448
rect 29536 158648 29592 159448
rect 30088 158648 30144 159448
rect 30732 158648 30788 159448
rect 31376 158648 31432 159448
rect 31928 158648 31984 159448
rect 32572 158648 32628 159448
rect 33216 158648 33272 159448
rect 33768 158648 33824 159448
rect 34412 158648 34468 159448
rect 35056 158648 35112 159448
rect 35608 158648 35664 159448
rect 36252 158648 36308 159448
rect 36896 158648 36952 159448
rect 37448 158648 37504 159448
rect 38092 158648 38148 159448
rect 38736 158648 38792 159448
rect 39380 158648 39436 159448
rect 39932 158648 39988 159448
rect 40576 158648 40632 159448
rect 41220 158648 41276 159448
rect 41772 158648 41828 159448
rect 42416 158648 42472 159448
rect 43060 158648 43116 159448
rect 43612 158648 43668 159448
rect 44256 158648 44312 159448
rect 44900 158648 44956 159448
rect 45452 158648 45508 159448
rect 46096 158648 46152 159448
rect 46740 158648 46796 159448
rect 47384 158648 47440 159448
rect 47936 158648 47992 159448
rect 48580 158648 48636 159448
rect 49224 158648 49280 159448
rect 49776 158648 49832 159448
rect 50420 158648 50476 159448
rect 51064 158648 51120 159448
rect 51616 158648 51672 159448
rect 52260 158648 52316 159448
rect 52904 158648 52960 159448
rect 53456 158648 53512 159448
rect 54100 158648 54156 159448
rect 54744 158648 54800 159448
rect 55296 158648 55352 159448
rect 55940 158648 55996 159448
rect 56584 158648 56640 159448
rect 57228 158648 57284 159448
rect 57780 158648 57836 159448
rect 58424 158648 58480 159448
rect 59068 158648 59124 159448
rect 59620 158648 59676 159448
rect 60264 158648 60320 159448
rect 60908 158648 60964 159448
rect 61460 158648 61516 159448
rect 62104 158648 62160 159448
rect 62748 158648 62804 159448
rect 63300 158648 63356 159448
rect 63944 158648 64000 159448
rect 64588 158648 64644 159448
rect 65140 158648 65196 159448
rect 65784 158648 65840 159448
rect 66428 158648 66484 159448
rect 67072 158648 67128 159448
rect 67624 158648 67680 159448
rect 68268 158648 68324 159448
rect 68912 158648 68968 159448
rect 69464 158648 69520 159448
rect 70108 158648 70164 159448
rect 70752 158648 70808 159448
rect 71304 158648 71360 159448
rect 71948 158648 72004 159448
rect 72592 158648 72648 159448
rect 73144 158648 73200 159448
rect 73788 158648 73844 159448
rect 74432 158648 74488 159448
rect 74984 158648 75040 159448
rect 75628 158648 75684 159448
rect 76272 158648 76328 159448
rect 76916 158648 76972 159448
rect 77468 158648 77524 159448
rect 78112 158648 78168 159448
rect 78756 158648 78812 159448
rect 79308 158648 79364 159448
rect 79952 158648 80008 159448
rect 80596 158648 80652 159448
rect 81148 158648 81204 159448
rect 81792 158648 81848 159448
rect 82436 158648 82492 159448
rect 82988 158648 83044 159448
rect 83632 158648 83688 159448
rect 84276 158648 84332 159448
rect 84920 158648 84976 159448
rect 85472 158648 85528 159448
rect 86116 158648 86172 159448
rect 86760 158648 86816 159448
rect 87312 158648 87368 159448
rect 87956 158648 88012 159448
rect 88600 158648 88656 159448
rect 89152 158648 89208 159448
rect 89796 158648 89852 159448
rect 90440 158648 90496 159448
rect 90992 158648 91048 159448
rect 91636 158648 91692 159448
rect 92280 158648 92336 159448
rect 92832 158648 92888 159448
rect 93476 158648 93532 159448
rect 94120 158648 94176 159448
rect 94764 158648 94820 159448
rect 95316 158648 95372 159448
rect 95960 158648 96016 159448
rect 96604 158648 96660 159448
rect 97156 158648 97212 159448
rect 97800 158648 97856 159448
rect 98444 158648 98500 159448
rect 98996 158648 99052 159448
rect 99640 158648 99696 159448
rect 100284 158648 100340 159448
rect 100836 158648 100892 159448
rect 101480 158648 101536 159448
rect 102124 158648 102180 159448
rect 102676 158648 102732 159448
rect 103320 158648 103376 159448
rect 103964 158648 104020 159448
rect 104608 158648 104664 159448
rect 105160 158648 105216 159448
rect 105804 158648 105860 159448
rect 106448 158648 106504 159448
rect 107000 158648 107056 159448
rect 107644 158648 107700 159448
rect 108288 158648 108344 159448
rect 108840 158648 108896 159448
rect 109484 158648 109540 159448
rect 110128 158648 110184 159448
rect 110680 158648 110736 159448
rect 111324 158648 111380 159448
rect 111968 158648 112024 159448
rect 112520 158648 112576 159448
rect 113164 158648 113220 159448
rect 113808 158648 113864 159448
rect 114452 158648 114508 159448
rect 115004 158648 115060 159448
rect 115648 158648 115704 159448
rect 116292 158648 116348 159448
rect 116844 158648 116900 159448
rect 117488 158648 117544 159448
rect 118132 158648 118188 159448
rect 118684 158648 118740 159448
rect 119328 158648 119384 159448
rect 119972 158648 120028 159448
rect 120524 158648 120580 159448
rect 121168 158648 121224 159448
rect 121812 158648 121868 159448
rect 122456 158648 122512 159448
rect 123008 158648 123064 159448
rect 123652 158648 123708 159448
rect 124296 158648 124352 159448
rect 124848 158648 124904 159448
rect 125492 158648 125548 159448
rect 126136 158648 126192 159448
rect 126688 158648 126744 159448
rect 127332 158648 127388 159448
rect 127976 158648 128032 159448
rect 128528 158648 128584 159448
rect 129172 158648 129228 159448
rect 129816 158648 129872 159448
rect 130368 158648 130424 159448
rect 131012 158648 131068 159448
rect 131656 158648 131712 159448
rect 132300 158648 132356 159448
rect 132852 158648 132908 159448
rect 133496 158648 133552 159448
rect 134140 158648 134196 159448
rect 134692 158648 134748 159448
rect 135336 158648 135392 159448
rect 135980 158648 136036 159448
rect 136532 158648 136588 159448
rect 137176 158648 137232 159448
rect 137820 158648 137876 159448
rect 138372 158648 138428 159448
rect 139016 158648 139072 159448
rect 139660 158648 139716 159448
rect 140212 158648 140268 159448
rect 140856 158648 140912 159448
rect 141500 158648 141556 159448
rect 142144 158648 142200 159448
rect 142696 158648 142752 159448
rect 143340 158648 143396 159448
rect 143984 158648 144040 159448
rect 144536 158648 144592 159448
rect 145180 158648 145236 159448
rect 145824 158648 145880 159448
rect 146376 158648 146432 159448
rect 147020 158648 147076 159448
rect 147664 158648 147720 159448
rect 148216 158648 148272 159448
rect 148860 158648 148916 159448
rect 149504 158648 149560 159448
rect 150056 158648 150112 159448
rect 150700 158648 150756 159448
rect 151344 158648 151400 159448
rect 151988 158648 152044 159448
rect 152540 158648 152596 159448
rect 153184 158648 153240 159448
rect 153828 158648 153884 159448
rect 154380 158648 154436 159448
rect 155024 158648 155080 159448
rect 155668 158648 155724 159448
rect 156220 158648 156276 159448
rect 156864 158648 156920 159448
rect 157508 158648 157564 159448
rect 158060 158648 158116 159448
rect 158704 158648 158760 159448
rect 159348 158648 159404 159448
<< obsm2 >>
rect 116 158592 500 158673
rect 668 158592 1144 158673
rect 1312 158592 1788 158673
rect 1956 158592 2340 158673
rect 2508 158592 2984 158673
rect 3152 158592 3628 158673
rect 3796 158592 4180 158673
rect 4348 158592 4824 158673
rect 4992 158592 5468 158673
rect 5636 158592 6020 158673
rect 6188 158592 6664 158673
rect 6832 158592 7308 158673
rect 7476 158592 7860 158673
rect 8028 158592 8504 158673
rect 8672 158592 9148 158673
rect 9316 158592 9792 158673
rect 9960 158592 10344 158673
rect 10512 158592 10988 158673
rect 11156 158592 11632 158673
rect 11800 158592 12184 158673
rect 12352 158592 12828 158673
rect 12996 158592 13472 158673
rect 13640 158592 14024 158673
rect 14192 158592 14668 158673
rect 14836 158592 15312 158673
rect 15480 158592 15864 158673
rect 16032 158592 16508 158673
rect 16676 158592 17152 158673
rect 17320 158592 17704 158673
rect 17872 158592 18348 158673
rect 18516 158592 18992 158673
rect 19160 158592 19636 158673
rect 19804 158592 20188 158673
rect 20356 158592 20832 158673
rect 21000 158592 21476 158673
rect 21644 158592 22028 158673
rect 22196 158592 22672 158673
rect 22840 158592 23316 158673
rect 23484 158592 23868 158673
rect 24036 158592 24512 158673
rect 24680 158592 25156 158673
rect 25324 158592 25708 158673
rect 25876 158592 26352 158673
rect 26520 158592 26996 158673
rect 27164 158592 27548 158673
rect 27716 158592 28192 158673
rect 28360 158592 28836 158673
rect 29004 158592 29480 158673
rect 29648 158592 30032 158673
rect 30200 158592 30676 158673
rect 30844 158592 31320 158673
rect 31488 158592 31872 158673
rect 32040 158592 32516 158673
rect 32684 158592 33160 158673
rect 33328 158592 33712 158673
rect 33880 158592 34356 158673
rect 34524 158592 35000 158673
rect 35168 158592 35552 158673
rect 35720 158592 36196 158673
rect 36364 158592 36840 158673
rect 37008 158592 37392 158673
rect 37560 158592 38036 158673
rect 38204 158592 38680 158673
rect 38848 158592 39324 158673
rect 39492 158592 39876 158673
rect 40044 158592 40520 158673
rect 40688 158592 41164 158673
rect 41332 158592 41716 158673
rect 41884 158592 42360 158673
rect 42528 158592 43004 158673
rect 43172 158592 43556 158673
rect 43724 158592 44200 158673
rect 44368 158592 44844 158673
rect 45012 158592 45396 158673
rect 45564 158592 46040 158673
rect 46208 158592 46684 158673
rect 46852 158592 47328 158673
rect 47496 158592 47880 158673
rect 48048 158592 48524 158673
rect 48692 158592 49168 158673
rect 49336 158592 49720 158673
rect 49888 158592 50364 158673
rect 50532 158592 51008 158673
rect 51176 158592 51560 158673
rect 51728 158592 52204 158673
rect 52372 158592 52848 158673
rect 53016 158592 53400 158673
rect 53568 158592 54044 158673
rect 54212 158592 54688 158673
rect 54856 158592 55240 158673
rect 55408 158592 55884 158673
rect 56052 158592 56528 158673
rect 56696 158592 57172 158673
rect 57340 158592 57724 158673
rect 57892 158592 58368 158673
rect 58536 158592 59012 158673
rect 59180 158592 59564 158673
rect 59732 158592 60208 158673
rect 60376 158592 60852 158673
rect 61020 158592 61404 158673
rect 61572 158592 62048 158673
rect 62216 158592 62692 158673
rect 62860 158592 63244 158673
rect 63412 158592 63888 158673
rect 64056 158592 64532 158673
rect 64700 158592 65084 158673
rect 65252 158592 65728 158673
rect 65896 158592 66372 158673
rect 66540 158592 67016 158673
rect 67184 158592 67568 158673
rect 67736 158592 68212 158673
rect 68380 158592 68856 158673
rect 69024 158592 69408 158673
rect 69576 158592 70052 158673
rect 70220 158592 70696 158673
rect 70864 158592 71248 158673
rect 71416 158592 71892 158673
rect 72060 158592 72536 158673
rect 72704 158592 73088 158673
rect 73256 158592 73732 158673
rect 73900 158592 74376 158673
rect 74544 158592 74928 158673
rect 75096 158592 75572 158673
rect 75740 158592 76216 158673
rect 76384 158592 76860 158673
rect 77028 158592 77412 158673
rect 77580 158592 78056 158673
rect 78224 158592 78700 158673
rect 78868 158592 79252 158673
rect 79420 158592 79896 158673
rect 80064 158592 80540 158673
rect 80708 158592 81092 158673
rect 81260 158592 81736 158673
rect 81904 158592 82380 158673
rect 82548 158592 82932 158673
rect 83100 158592 83576 158673
rect 83744 158592 84220 158673
rect 84388 158592 84864 158673
rect 85032 158592 85416 158673
rect 85584 158592 86060 158673
rect 86228 158592 86704 158673
rect 86872 158592 87256 158673
rect 87424 158592 87900 158673
rect 88068 158592 88544 158673
rect 88712 158592 89096 158673
rect 89264 158592 89740 158673
rect 89908 158592 90384 158673
rect 90552 158592 90936 158673
rect 91104 158592 91580 158673
rect 91748 158592 92224 158673
rect 92392 158592 92776 158673
rect 92944 158592 93420 158673
rect 93588 158592 94064 158673
rect 94232 158592 94708 158673
rect 94876 158592 95260 158673
rect 95428 158592 95904 158673
rect 96072 158592 96548 158673
rect 96716 158592 97100 158673
rect 97268 158592 97744 158673
rect 97912 158592 98388 158673
rect 98556 158592 98940 158673
rect 99108 158592 99584 158673
rect 99752 158592 100228 158673
rect 100396 158592 100780 158673
rect 100948 158592 101424 158673
rect 101592 158592 102068 158673
rect 102236 158592 102620 158673
rect 102788 158592 103264 158673
rect 103432 158592 103908 158673
rect 104076 158592 104552 158673
rect 104720 158592 105104 158673
rect 105272 158592 105748 158673
rect 105916 158592 106392 158673
rect 106560 158592 106944 158673
rect 107112 158592 107588 158673
rect 107756 158592 108232 158673
rect 108400 158592 108784 158673
rect 108952 158592 109428 158673
rect 109596 158592 110072 158673
rect 110240 158592 110624 158673
rect 110792 158592 111268 158673
rect 111436 158592 111912 158673
rect 112080 158592 112464 158673
rect 112632 158592 113108 158673
rect 113276 158592 113752 158673
rect 113920 158592 114396 158673
rect 114564 158592 114948 158673
rect 115116 158592 115592 158673
rect 115760 158592 116236 158673
rect 116404 158592 116788 158673
rect 116956 158592 117432 158673
rect 117600 158592 118076 158673
rect 118244 158592 118628 158673
rect 118796 158592 119272 158673
rect 119440 158592 119916 158673
rect 120084 158592 120468 158673
rect 120636 158592 121112 158673
rect 121280 158592 121756 158673
rect 121924 158592 122400 158673
rect 122568 158592 122952 158673
rect 123120 158592 123596 158673
rect 123764 158592 124240 158673
rect 124408 158592 124792 158673
rect 124960 158592 125436 158673
rect 125604 158592 126080 158673
rect 126248 158592 126632 158673
rect 126800 158592 127276 158673
rect 127444 158592 127920 158673
rect 128088 158592 128472 158673
rect 128640 158592 129116 158673
rect 129284 158592 129760 158673
rect 129928 158592 130312 158673
rect 130480 158592 130956 158673
rect 131124 158592 131600 158673
rect 131768 158592 132244 158673
rect 132412 158592 132796 158673
rect 132964 158592 133440 158673
rect 133608 158592 134084 158673
rect 134252 158592 134636 158673
rect 134804 158592 135280 158673
rect 135448 158592 135924 158673
rect 136092 158592 136476 158673
rect 136644 158592 137120 158673
rect 137288 158592 137764 158673
rect 137932 158592 138316 158673
rect 138484 158592 138960 158673
rect 139128 158592 139604 158673
rect 139772 158592 140156 158673
rect 140324 158592 140800 158673
rect 140968 158592 141444 158673
rect 141612 158592 142088 158673
rect 142256 158592 142640 158673
rect 142808 158592 143284 158673
rect 143452 158592 143928 158673
rect 144096 158592 144480 158673
rect 144648 158592 145124 158673
rect 145292 158592 145768 158673
rect 145936 158592 146320 158673
rect 146488 158592 146964 158673
rect 147132 158592 147608 158673
rect 147776 158592 148160 158673
rect 148328 158592 148804 158673
rect 148972 158592 149448 158673
rect 149616 158592 150000 158673
rect 150168 158592 150644 158673
rect 150812 158592 151288 158673
rect 151456 158592 151932 158673
rect 152100 158592 152484 158673
rect 152652 158592 153128 158673
rect 153296 158592 153772 158673
rect 153940 158592 154324 158673
rect 154492 158592 154968 158673
rect 155136 158592 155612 158673
rect 155780 158592 156164 158673
rect 156332 158592 156808 158673
rect 156976 158592 157452 158673
rect 157620 158592 158004 158673
rect 158172 158592 158648 158673
rect 158816 158592 159292 158673
rect 6 23 159402 158592
<< metal3 >>
rect 158910 158576 159710 158696
rect 158910 157352 159710 157472
rect 158910 156128 159710 156248
rect 158910 154904 159710 155024
rect 158910 153680 159710 153800
rect 158910 152456 159710 152576
rect 158910 151232 159710 151352
rect 158910 150008 159710 150128
rect 158910 148784 159710 148904
rect 158910 147560 159710 147680
rect 158910 146336 159710 146456
rect 158910 145112 159710 145232
rect 158910 143888 159710 144008
rect 158910 142664 159710 142784
rect 158910 141440 159710 141560
rect 158910 140216 159710 140336
rect 158910 138992 159710 139112
rect 158910 137768 159710 137888
rect 158910 136544 159710 136664
rect 158910 135320 159710 135440
rect 158910 134096 159710 134216
rect 158910 132736 159710 132856
rect 158910 131512 159710 131632
rect 158910 130288 159710 130408
rect 158910 129064 159710 129184
rect 158910 127840 159710 127960
rect 158910 126616 159710 126736
rect 158910 125392 159710 125512
rect 158910 124168 159710 124288
rect 158910 122944 159710 123064
rect 158910 121720 159710 121840
rect 158910 120496 159710 120616
rect 158910 119272 159710 119392
rect 158910 118048 159710 118168
rect 158910 116824 159710 116944
rect 158910 115600 159710 115720
rect 158910 114376 159710 114496
rect 158910 113152 159710 113272
rect 158910 111928 159710 112048
rect 158910 110704 159710 110824
rect 158910 109480 159710 109600
rect 158910 108256 159710 108376
rect 158910 107032 159710 107152
rect 158910 105672 159710 105792
rect 158910 104448 159710 104568
rect 158910 103224 159710 103344
rect 158910 102000 159710 102120
rect 158910 100776 159710 100896
rect 158910 99552 159710 99672
rect 158910 98328 159710 98448
rect 158910 97104 159710 97224
rect 158910 95880 159710 96000
rect 158910 94656 159710 94776
rect 158910 93432 159710 93552
rect 158910 92208 159710 92328
rect 158910 90984 159710 91104
rect 158910 89760 159710 89880
rect 158910 88536 159710 88656
rect 158910 87312 159710 87432
rect 158910 86088 159710 86208
rect 158910 84864 159710 84984
rect 158910 83640 159710 83760
rect 158910 82416 159710 82536
rect 158910 81192 159710 81312
rect 158910 79968 159710 80088
rect 158910 78608 159710 78728
rect 158910 77384 159710 77504
rect 158910 76160 159710 76280
rect 158910 74936 159710 75056
rect 158910 73712 159710 73832
rect 158910 72488 159710 72608
rect 158910 71264 159710 71384
rect 158910 70040 159710 70160
rect 158910 68816 159710 68936
rect 158910 67592 159710 67712
rect 158910 66368 159710 66488
rect 158910 65144 159710 65264
rect 158910 63920 159710 64040
rect 158910 62696 159710 62816
rect 158910 61472 159710 61592
rect 158910 60248 159710 60368
rect 158910 59024 159710 59144
rect 158910 57800 159710 57920
rect 158910 56576 159710 56696
rect 158910 55352 159710 55472
rect 158910 54128 159710 54248
rect 158910 52768 159710 52888
rect 158910 51544 159710 51664
rect 158910 50320 159710 50440
rect 158910 49096 159710 49216
rect 158910 47872 159710 47992
rect 158910 46648 159710 46768
rect 158910 45424 159710 45544
rect 158910 44200 159710 44320
rect 158910 42976 159710 43096
rect 158910 41752 159710 41872
rect 158910 40528 159710 40648
rect 158910 39304 159710 39424
rect 158910 38080 159710 38200
rect 158910 36856 159710 36976
rect 158910 35632 159710 35752
rect 158910 34408 159710 34528
rect 158910 33184 159710 33304
rect 158910 31960 159710 32080
rect 158910 30736 159710 30856
rect 158910 29512 159710 29632
rect 158910 28288 159710 28408
rect 158910 27064 159710 27184
rect 158910 25704 159710 25824
rect 158910 24480 159710 24600
rect 158910 23256 159710 23376
rect 158910 22032 159710 22152
rect 158910 20808 159710 20928
rect 158910 19584 159710 19704
rect 158910 18360 159710 18480
rect 158910 17136 159710 17256
rect 158910 15912 159710 16032
rect 158910 14688 159710 14808
rect 158910 13464 159710 13584
rect 158910 12240 159710 12360
rect 158910 11016 159710 11136
rect 158910 9792 159710 9912
rect 158910 8568 159710 8688
rect 158910 7344 159710 7464
rect 158910 6120 159710 6240
rect 158910 4896 159710 5016
rect 158910 3672 159710 3792
rect 158910 2448 159710 2568
rect 158910 1224 159710 1344
rect 158910 0 159710 120
<< obsm3 >>
rect 1379 158496 158830 158669
rect 1379 157552 159041 158496
rect 1379 157272 158830 157552
rect 1379 156328 159041 157272
rect 1379 156048 158830 156328
rect 1379 155104 159041 156048
rect 1379 154824 158830 155104
rect 1379 153880 159041 154824
rect 1379 153600 158830 153880
rect 1379 152656 159041 153600
rect 1379 152376 158830 152656
rect 1379 151432 159041 152376
rect 1379 151152 158830 151432
rect 1379 150208 159041 151152
rect 1379 149928 158830 150208
rect 1379 148984 159041 149928
rect 1379 148704 158830 148984
rect 1379 147760 159041 148704
rect 1379 147480 158830 147760
rect 1379 146536 159041 147480
rect 1379 146256 158830 146536
rect 1379 145312 159041 146256
rect 1379 145032 158830 145312
rect 1379 144088 159041 145032
rect 1379 143808 158830 144088
rect 1379 142864 159041 143808
rect 1379 142584 158830 142864
rect 1379 141640 159041 142584
rect 1379 141360 158830 141640
rect 1379 140416 159041 141360
rect 1379 140136 158830 140416
rect 1379 139192 159041 140136
rect 1379 138912 158830 139192
rect 1379 137968 159041 138912
rect 1379 137688 158830 137968
rect 1379 136744 159041 137688
rect 1379 136464 158830 136744
rect 1379 135520 159041 136464
rect 1379 135240 158830 135520
rect 1379 134296 159041 135240
rect 1379 134016 158830 134296
rect 1379 132936 159041 134016
rect 1379 132656 158830 132936
rect 1379 131712 159041 132656
rect 1379 131432 158830 131712
rect 1379 130488 159041 131432
rect 1379 130208 158830 130488
rect 1379 129264 159041 130208
rect 1379 128984 158830 129264
rect 1379 128040 159041 128984
rect 1379 127760 158830 128040
rect 1379 126816 159041 127760
rect 1379 126536 158830 126816
rect 1379 125592 159041 126536
rect 1379 125312 158830 125592
rect 1379 124368 159041 125312
rect 1379 124088 158830 124368
rect 1379 123144 159041 124088
rect 1379 122864 158830 123144
rect 1379 121920 159041 122864
rect 1379 121640 158830 121920
rect 1379 120696 159041 121640
rect 1379 120416 158830 120696
rect 1379 119472 159041 120416
rect 1379 119192 158830 119472
rect 1379 118248 159041 119192
rect 1379 117968 158830 118248
rect 1379 117024 159041 117968
rect 1379 116744 158830 117024
rect 1379 115800 159041 116744
rect 1379 115520 158830 115800
rect 1379 114576 159041 115520
rect 1379 114296 158830 114576
rect 1379 113352 159041 114296
rect 1379 113072 158830 113352
rect 1379 112128 159041 113072
rect 1379 111848 158830 112128
rect 1379 110904 159041 111848
rect 1379 110624 158830 110904
rect 1379 109680 159041 110624
rect 1379 109400 158830 109680
rect 1379 108456 159041 109400
rect 1379 108176 158830 108456
rect 1379 107232 159041 108176
rect 1379 106952 158830 107232
rect 1379 105872 159041 106952
rect 1379 105592 158830 105872
rect 1379 104648 159041 105592
rect 1379 104368 158830 104648
rect 1379 103424 159041 104368
rect 1379 103144 158830 103424
rect 1379 102200 159041 103144
rect 1379 101920 158830 102200
rect 1379 100976 159041 101920
rect 1379 100696 158830 100976
rect 1379 99752 159041 100696
rect 1379 99472 158830 99752
rect 1379 98528 159041 99472
rect 1379 98248 158830 98528
rect 1379 97304 159041 98248
rect 1379 97024 158830 97304
rect 1379 96080 159041 97024
rect 1379 95800 158830 96080
rect 1379 94856 159041 95800
rect 1379 94576 158830 94856
rect 1379 93632 159041 94576
rect 1379 93352 158830 93632
rect 1379 92408 159041 93352
rect 1379 92128 158830 92408
rect 1379 91184 159041 92128
rect 1379 90904 158830 91184
rect 1379 89960 159041 90904
rect 1379 89680 158830 89960
rect 1379 88736 159041 89680
rect 1379 88456 158830 88736
rect 1379 87512 159041 88456
rect 1379 87232 158830 87512
rect 1379 86288 159041 87232
rect 1379 86008 158830 86288
rect 1379 85064 159041 86008
rect 1379 84784 158830 85064
rect 1379 83840 159041 84784
rect 1379 83560 158830 83840
rect 1379 82616 159041 83560
rect 1379 82336 158830 82616
rect 1379 81392 159041 82336
rect 1379 81112 158830 81392
rect 1379 80168 159041 81112
rect 1379 79888 158830 80168
rect 1379 78808 159041 79888
rect 1379 78528 158830 78808
rect 1379 77584 159041 78528
rect 1379 77304 158830 77584
rect 1379 76360 159041 77304
rect 1379 76080 158830 76360
rect 1379 75136 159041 76080
rect 1379 74856 158830 75136
rect 1379 73912 159041 74856
rect 1379 73632 158830 73912
rect 1379 72688 159041 73632
rect 1379 72408 158830 72688
rect 1379 71464 159041 72408
rect 1379 71184 158830 71464
rect 1379 70240 159041 71184
rect 1379 69960 158830 70240
rect 1379 69016 159041 69960
rect 1379 68736 158830 69016
rect 1379 67792 159041 68736
rect 1379 67512 158830 67792
rect 1379 66568 159041 67512
rect 1379 66288 158830 66568
rect 1379 65344 159041 66288
rect 1379 65064 158830 65344
rect 1379 64120 159041 65064
rect 1379 63840 158830 64120
rect 1379 62896 159041 63840
rect 1379 62616 158830 62896
rect 1379 61672 159041 62616
rect 1379 61392 158830 61672
rect 1379 60448 159041 61392
rect 1379 60168 158830 60448
rect 1379 59224 159041 60168
rect 1379 58944 158830 59224
rect 1379 58000 159041 58944
rect 1379 57720 158830 58000
rect 1379 56776 159041 57720
rect 1379 56496 158830 56776
rect 1379 55552 159041 56496
rect 1379 55272 158830 55552
rect 1379 54328 159041 55272
rect 1379 54048 158830 54328
rect 1379 52968 159041 54048
rect 1379 52688 158830 52968
rect 1379 51744 159041 52688
rect 1379 51464 158830 51744
rect 1379 50520 159041 51464
rect 1379 50240 158830 50520
rect 1379 49296 159041 50240
rect 1379 49016 158830 49296
rect 1379 48072 159041 49016
rect 1379 47792 158830 48072
rect 1379 46848 159041 47792
rect 1379 46568 158830 46848
rect 1379 45624 159041 46568
rect 1379 45344 158830 45624
rect 1379 44400 159041 45344
rect 1379 44120 158830 44400
rect 1379 43176 159041 44120
rect 1379 42896 158830 43176
rect 1379 41952 159041 42896
rect 1379 41672 158830 41952
rect 1379 40728 159041 41672
rect 1379 40448 158830 40728
rect 1379 39504 159041 40448
rect 1379 39224 158830 39504
rect 1379 38280 159041 39224
rect 1379 38000 158830 38280
rect 1379 37056 159041 38000
rect 1379 36776 158830 37056
rect 1379 35832 159041 36776
rect 1379 35552 158830 35832
rect 1379 34608 159041 35552
rect 1379 34328 158830 34608
rect 1379 33384 159041 34328
rect 1379 33104 158830 33384
rect 1379 32160 159041 33104
rect 1379 31880 158830 32160
rect 1379 30936 159041 31880
rect 1379 30656 158830 30936
rect 1379 29712 159041 30656
rect 1379 29432 158830 29712
rect 1379 28488 159041 29432
rect 1379 28208 158830 28488
rect 1379 27264 159041 28208
rect 1379 26984 158830 27264
rect 1379 25904 159041 26984
rect 1379 25624 158830 25904
rect 1379 24680 159041 25624
rect 1379 24400 158830 24680
rect 1379 23456 159041 24400
rect 1379 23176 158830 23456
rect 1379 22232 159041 23176
rect 1379 21952 158830 22232
rect 1379 21008 159041 21952
rect 1379 20728 158830 21008
rect 1379 19784 159041 20728
rect 1379 19504 158830 19784
rect 1379 18560 159041 19504
rect 1379 18280 158830 18560
rect 1379 17336 159041 18280
rect 1379 17056 158830 17336
rect 1379 16112 159041 17056
rect 1379 15832 158830 16112
rect 1379 14888 159041 15832
rect 1379 14608 158830 14888
rect 1379 13664 159041 14608
rect 1379 13384 158830 13664
rect 1379 12440 159041 13384
rect 1379 12160 158830 12440
rect 1379 11216 159041 12160
rect 1379 10936 158830 11216
rect 1379 9992 159041 10936
rect 1379 9712 158830 9992
rect 1379 8768 159041 9712
rect 1379 8488 158830 8768
rect 1379 7544 159041 8488
rect 1379 7264 158830 7544
rect 1379 6320 159041 7264
rect 1379 6040 158830 6320
rect 1379 5096 159041 6040
rect 1379 4816 158830 5096
rect 1379 3872 159041 4816
rect 1379 3592 158830 3872
rect 1379 2648 159041 3592
rect 1379 2368 158830 2648
rect 1379 1424 159041 2368
rect 1379 1144 158830 1424
rect 1379 200 159041 1144
rect 1379 27 158830 200
<< metal4 >>
rect 3918 1576 4238 157256
rect 4578 1624 4898 157208
rect 5238 1624 5558 157208
rect 5898 1624 6218 157208
rect 19278 1576 19598 157256
rect 19938 1624 20258 157208
rect 20598 1624 20918 157208
rect 21258 1624 21578 157208
rect 34638 1576 34958 157256
rect 35298 1624 35618 157208
rect 35958 1624 36278 157208
rect 36618 1624 36938 157208
rect 49998 1576 50318 157256
rect 50658 1624 50978 157208
rect 51318 1624 51638 157208
rect 51978 1624 52298 157208
rect 65358 1576 65678 157256
rect 66018 1624 66338 157208
rect 66678 1624 66998 157208
rect 67338 1624 67658 157208
rect 80718 1576 81038 157256
rect 81378 1624 81698 157208
rect 82038 1624 82358 157208
rect 82698 1624 83018 157208
rect 96078 1576 96398 157256
rect 96738 1624 97058 157208
rect 97398 1624 97718 157208
rect 98058 1624 98378 157208
rect 111438 1576 111758 157256
rect 112098 1624 112418 157208
rect 112758 1624 113078 157208
rect 113418 1624 113738 157208
rect 126798 1576 127118 157256
rect 127458 1624 127778 157208
rect 128118 1624 128438 157208
rect 128778 1624 129098 157208
rect 142158 1576 142478 157256
rect 142818 1624 143138 157208
rect 143478 1624 143798 157208
rect 144138 1624 144458 157208
rect 157518 1576 157838 157256
<< obsm4 >>
rect 2897 4107 3838 157309
rect 4318 157288 19198 157309
rect 4318 4107 4498 157288
rect 4978 4107 5158 157288
rect 5638 4107 5818 157288
rect 6298 4107 19198 157288
rect 19678 157288 34558 157309
rect 19678 4107 19858 157288
rect 20338 4107 20518 157288
rect 20998 4107 21178 157288
rect 21658 4107 34558 157288
rect 35038 157288 49918 157309
rect 35038 4107 35218 157288
rect 35698 4107 35878 157288
rect 36358 4107 36538 157288
rect 37018 4107 49918 157288
rect 50398 157288 65278 157309
rect 50398 4107 50578 157288
rect 51058 4107 51238 157288
rect 51718 4107 51898 157288
rect 52378 4107 65278 157288
rect 65758 157288 80638 157309
rect 65758 4107 65938 157288
rect 66418 4107 66598 157288
rect 67078 4107 67258 157288
rect 67738 4107 80638 157288
rect 81118 157288 95998 157309
rect 81118 4107 81298 157288
rect 81778 4107 81958 157288
rect 82438 4107 82618 157288
rect 83098 4107 95998 157288
rect 96478 157288 111358 157309
rect 96478 4107 96658 157288
rect 97138 4107 97318 157288
rect 97798 4107 97978 157288
rect 98458 4107 111358 157288
rect 111838 157288 126718 157309
rect 111838 4107 112018 157288
rect 112498 4107 112678 157288
rect 113158 4107 113338 157288
rect 113818 4107 126718 157288
rect 127198 157288 142078 157309
rect 127198 4107 127378 157288
rect 127858 4107 128038 157288
rect 128518 4107 128698 157288
rect 129178 4107 142078 157288
rect 142558 157288 157339 157309
rect 142558 4107 142738 157288
rect 143218 4107 143398 157288
rect 143878 4107 144058 157288
rect 144538 4107 157339 157288
<< labels >>
rlabel metal2 s 159348 158648 159404 159448 6 clk
port 1 nsew signal input
rlabel metal2 s 4 158648 60 159448 6 m_in[0]
port 2 nsew signal input
rlabel metal2 s 61460 158648 61516 159448 6 m_in[100]
port 3 nsew signal input
rlabel metal2 s 62104 158648 62160 159448 6 m_in[101]
port 4 nsew signal input
rlabel metal2 s 62748 158648 62804 159448 6 m_in[102]
port 5 nsew signal input
rlabel metal2 s 63300 158648 63356 159448 6 m_in[103]
port 6 nsew signal input
rlabel metal2 s 63944 158648 64000 159448 6 m_in[104]
port 7 nsew signal input
rlabel metal2 s 64588 158648 64644 159448 6 m_in[105]
port 8 nsew signal input
rlabel metal2 s 65140 158648 65196 159448 6 m_in[106]
port 9 nsew signal input
rlabel metal2 s 65784 158648 65840 159448 6 m_in[107]
port 10 nsew signal input
rlabel metal2 s 66428 158648 66484 159448 6 m_in[108]
port 11 nsew signal input
rlabel metal2 s 67072 158648 67128 159448 6 m_in[109]
port 12 nsew signal input
rlabel metal2 s 6076 158648 6132 159448 6 m_in[10]
port 13 nsew signal input
rlabel metal2 s 67624 158648 67680 159448 6 m_in[110]
port 14 nsew signal input
rlabel metal2 s 68268 158648 68324 159448 6 m_in[111]
port 15 nsew signal input
rlabel metal2 s 68912 158648 68968 159448 6 m_in[112]
port 16 nsew signal input
rlabel metal2 s 69464 158648 69520 159448 6 m_in[113]
port 17 nsew signal input
rlabel metal2 s 70108 158648 70164 159448 6 m_in[114]
port 18 nsew signal input
rlabel metal2 s 70752 158648 70808 159448 6 m_in[115]
port 19 nsew signal input
rlabel metal2 s 71304 158648 71360 159448 6 m_in[116]
port 20 nsew signal input
rlabel metal2 s 71948 158648 72004 159448 6 m_in[117]
port 21 nsew signal input
rlabel metal2 s 72592 158648 72648 159448 6 m_in[118]
port 22 nsew signal input
rlabel metal2 s 73144 158648 73200 159448 6 m_in[119]
port 23 nsew signal input
rlabel metal2 s 6720 158648 6776 159448 6 m_in[11]
port 24 nsew signal input
rlabel metal2 s 73788 158648 73844 159448 6 m_in[120]
port 25 nsew signal input
rlabel metal2 s 74432 158648 74488 159448 6 m_in[121]
port 26 nsew signal input
rlabel metal2 s 74984 158648 75040 159448 6 m_in[122]
port 27 nsew signal input
rlabel metal2 s 75628 158648 75684 159448 6 m_in[123]
port 28 nsew signal input
rlabel metal2 s 76272 158648 76328 159448 6 m_in[124]
port 29 nsew signal input
rlabel metal2 s 76916 158648 76972 159448 6 m_in[125]
port 30 nsew signal input
rlabel metal2 s 77468 158648 77524 159448 6 m_in[126]
port 31 nsew signal input
rlabel metal2 s 78112 158648 78168 159448 6 m_in[127]
port 32 nsew signal input
rlabel metal2 s 78756 158648 78812 159448 6 m_in[128]
port 33 nsew signal input
rlabel metal2 s 79308 158648 79364 159448 6 m_in[129]
port 34 nsew signal input
rlabel metal2 s 7364 158648 7420 159448 6 m_in[12]
port 35 nsew signal input
rlabel metal2 s 79952 158648 80008 159448 6 m_in[130]
port 36 nsew signal input
rlabel metal2 s 80596 158648 80652 159448 6 m_in[131]
port 37 nsew signal input
rlabel metal2 s 81148 158648 81204 159448 6 m_in[132]
port 38 nsew signal input
rlabel metal2 s 81792 158648 81848 159448 6 m_in[133]
port 39 nsew signal input
rlabel metal2 s 82436 158648 82492 159448 6 m_in[134]
port 40 nsew signal input
rlabel metal2 s 82988 158648 83044 159448 6 m_in[135]
port 41 nsew signal input
rlabel metal2 s 83632 158648 83688 159448 6 m_in[136]
port 42 nsew signal input
rlabel metal2 s 84276 158648 84332 159448 6 m_in[137]
port 43 nsew signal input
rlabel metal2 s 84920 158648 84976 159448 6 m_in[138]
port 44 nsew signal input
rlabel metal2 s 85472 158648 85528 159448 6 m_in[139]
port 45 nsew signal input
rlabel metal2 s 7916 158648 7972 159448 6 m_in[13]
port 46 nsew signal input
rlabel metal2 s 86116 158648 86172 159448 6 m_in[140]
port 47 nsew signal input
rlabel metal2 s 86760 158648 86816 159448 6 m_in[141]
port 48 nsew signal input
rlabel metal2 s 87312 158648 87368 159448 6 m_in[142]
port 49 nsew signal input
rlabel metal2 s 87956 158648 88012 159448 6 m_in[143]
port 50 nsew signal input
rlabel metal2 s 88600 158648 88656 159448 6 m_in[144]
port 51 nsew signal input
rlabel metal2 s 89152 158648 89208 159448 6 m_in[145]
port 52 nsew signal input
rlabel metal2 s 89796 158648 89852 159448 6 m_in[146]
port 53 nsew signal input
rlabel metal2 s 90440 158648 90496 159448 6 m_in[147]
port 54 nsew signal input
rlabel metal2 s 90992 158648 91048 159448 6 m_in[148]
port 55 nsew signal input
rlabel metal2 s 91636 158648 91692 159448 6 m_in[149]
port 56 nsew signal input
rlabel metal2 s 8560 158648 8616 159448 6 m_in[14]
port 57 nsew signal input
rlabel metal2 s 92280 158648 92336 159448 6 m_in[150]
port 58 nsew signal input
rlabel metal2 s 92832 158648 92888 159448 6 m_in[151]
port 59 nsew signal input
rlabel metal2 s 93476 158648 93532 159448 6 m_in[152]
port 60 nsew signal input
rlabel metal2 s 94120 158648 94176 159448 6 m_in[153]
port 61 nsew signal input
rlabel metal2 s 94764 158648 94820 159448 6 m_in[154]
port 62 nsew signal input
rlabel metal2 s 95316 158648 95372 159448 6 m_in[155]
port 63 nsew signal input
rlabel metal2 s 95960 158648 96016 159448 6 m_in[156]
port 64 nsew signal input
rlabel metal2 s 96604 158648 96660 159448 6 m_in[157]
port 65 nsew signal input
rlabel metal2 s 97156 158648 97212 159448 6 m_in[158]
port 66 nsew signal input
rlabel metal2 s 97800 158648 97856 159448 6 m_in[159]
port 67 nsew signal input
rlabel metal2 s 9204 158648 9260 159448 6 m_in[15]
port 68 nsew signal input
rlabel metal2 s 98444 158648 98500 159448 6 m_in[160]
port 69 nsew signal input
rlabel metal2 s 98996 158648 99052 159448 6 m_in[161]
port 70 nsew signal input
rlabel metal2 s 99640 158648 99696 159448 6 m_in[162]
port 71 nsew signal input
rlabel metal2 s 100284 158648 100340 159448 6 m_in[163]
port 72 nsew signal input
rlabel metal2 s 100836 158648 100892 159448 6 m_in[164]
port 73 nsew signal input
rlabel metal2 s 101480 158648 101536 159448 6 m_in[165]
port 74 nsew signal input
rlabel metal2 s 102124 158648 102180 159448 6 m_in[166]
port 75 nsew signal input
rlabel metal2 s 102676 158648 102732 159448 6 m_in[167]
port 76 nsew signal input
rlabel metal2 s 103320 158648 103376 159448 6 m_in[168]
port 77 nsew signal input
rlabel metal2 s 103964 158648 104020 159448 6 m_in[169]
port 78 nsew signal input
rlabel metal2 s 9848 158648 9904 159448 6 m_in[16]
port 79 nsew signal input
rlabel metal2 s 104608 158648 104664 159448 6 m_in[170]
port 80 nsew signal input
rlabel metal2 s 105160 158648 105216 159448 6 m_in[171]
port 81 nsew signal input
rlabel metal2 s 105804 158648 105860 159448 6 m_in[172]
port 82 nsew signal input
rlabel metal2 s 106448 158648 106504 159448 6 m_in[173]
port 83 nsew signal input
rlabel metal2 s 107000 158648 107056 159448 6 m_in[174]
port 84 nsew signal input
rlabel metal2 s 107644 158648 107700 159448 6 m_in[175]
port 85 nsew signal input
rlabel metal2 s 108288 158648 108344 159448 6 m_in[176]
port 86 nsew signal input
rlabel metal2 s 108840 158648 108896 159448 6 m_in[177]
port 87 nsew signal input
rlabel metal2 s 109484 158648 109540 159448 6 m_in[178]
port 88 nsew signal input
rlabel metal2 s 110128 158648 110184 159448 6 m_in[179]
port 89 nsew signal input
rlabel metal2 s 10400 158648 10456 159448 6 m_in[17]
port 90 nsew signal input
rlabel metal2 s 110680 158648 110736 159448 6 m_in[180]
port 91 nsew signal input
rlabel metal2 s 111324 158648 111380 159448 6 m_in[181]
port 92 nsew signal input
rlabel metal2 s 111968 158648 112024 159448 6 m_in[182]
port 93 nsew signal input
rlabel metal2 s 112520 158648 112576 159448 6 m_in[183]
port 94 nsew signal input
rlabel metal2 s 113164 158648 113220 159448 6 m_in[184]
port 95 nsew signal input
rlabel metal2 s 113808 158648 113864 159448 6 m_in[185]
port 96 nsew signal input
rlabel metal2 s 114452 158648 114508 159448 6 m_in[186]
port 97 nsew signal input
rlabel metal2 s 115004 158648 115060 159448 6 m_in[187]
port 98 nsew signal input
rlabel metal2 s 115648 158648 115704 159448 6 m_in[188]
port 99 nsew signal input
rlabel metal2 s 116292 158648 116348 159448 6 m_in[189]
port 100 nsew signal input
rlabel metal2 s 11044 158648 11100 159448 6 m_in[18]
port 101 nsew signal input
rlabel metal2 s 116844 158648 116900 159448 6 m_in[190]
port 102 nsew signal input
rlabel metal2 s 117488 158648 117544 159448 6 m_in[191]
port 103 nsew signal input
rlabel metal2 s 118132 158648 118188 159448 6 m_in[192]
port 104 nsew signal input
rlabel metal2 s 118684 158648 118740 159448 6 m_in[193]
port 105 nsew signal input
rlabel metal2 s 119328 158648 119384 159448 6 m_in[194]
port 106 nsew signal input
rlabel metal2 s 119972 158648 120028 159448 6 m_in[195]
port 107 nsew signal input
rlabel metal2 s 120524 158648 120580 159448 6 m_in[196]
port 108 nsew signal input
rlabel metal2 s 121168 158648 121224 159448 6 m_in[197]
port 109 nsew signal input
rlabel metal2 s 121812 158648 121868 159448 6 m_in[198]
port 110 nsew signal input
rlabel metal2 s 122456 158648 122512 159448 6 m_in[199]
port 111 nsew signal input
rlabel metal2 s 11688 158648 11744 159448 6 m_in[19]
port 112 nsew signal input
rlabel metal2 s 556 158648 612 159448 6 m_in[1]
port 113 nsew signal input
rlabel metal2 s 123008 158648 123064 159448 6 m_in[200]
port 114 nsew signal input
rlabel metal2 s 123652 158648 123708 159448 6 m_in[201]
port 115 nsew signal input
rlabel metal2 s 124296 158648 124352 159448 6 m_in[202]
port 116 nsew signal input
rlabel metal2 s 124848 158648 124904 159448 6 m_in[203]
port 117 nsew signal input
rlabel metal2 s 125492 158648 125548 159448 6 m_in[204]
port 118 nsew signal input
rlabel metal2 s 126136 158648 126192 159448 6 m_in[205]
port 119 nsew signal input
rlabel metal2 s 126688 158648 126744 159448 6 m_in[206]
port 120 nsew signal input
rlabel metal2 s 127332 158648 127388 159448 6 m_in[207]
port 121 nsew signal input
rlabel metal2 s 127976 158648 128032 159448 6 m_in[208]
port 122 nsew signal input
rlabel metal2 s 128528 158648 128584 159448 6 m_in[209]
port 123 nsew signal input
rlabel metal2 s 12240 158648 12296 159448 6 m_in[20]
port 124 nsew signal input
rlabel metal2 s 129172 158648 129228 159448 6 m_in[210]
port 125 nsew signal input
rlabel metal2 s 129816 158648 129872 159448 6 m_in[211]
port 126 nsew signal input
rlabel metal2 s 130368 158648 130424 159448 6 m_in[212]
port 127 nsew signal input
rlabel metal2 s 131012 158648 131068 159448 6 m_in[213]
port 128 nsew signal input
rlabel metal2 s 131656 158648 131712 159448 6 m_in[214]
port 129 nsew signal input
rlabel metal2 s 132300 158648 132356 159448 6 m_in[215]
port 130 nsew signal input
rlabel metal2 s 132852 158648 132908 159448 6 m_in[216]
port 131 nsew signal input
rlabel metal2 s 133496 158648 133552 159448 6 m_in[217]
port 132 nsew signal input
rlabel metal2 s 134140 158648 134196 159448 6 m_in[218]
port 133 nsew signal input
rlabel metal2 s 134692 158648 134748 159448 6 m_in[219]
port 134 nsew signal input
rlabel metal2 s 12884 158648 12940 159448 6 m_in[21]
port 135 nsew signal input
rlabel metal2 s 135336 158648 135392 159448 6 m_in[220]
port 136 nsew signal input
rlabel metal2 s 135980 158648 136036 159448 6 m_in[221]
port 137 nsew signal input
rlabel metal2 s 136532 158648 136588 159448 6 m_in[222]
port 138 nsew signal input
rlabel metal2 s 137176 158648 137232 159448 6 m_in[223]
port 139 nsew signal input
rlabel metal2 s 137820 158648 137876 159448 6 m_in[224]
port 140 nsew signal input
rlabel metal2 s 138372 158648 138428 159448 6 m_in[225]
port 141 nsew signal input
rlabel metal2 s 139016 158648 139072 159448 6 m_in[226]
port 142 nsew signal input
rlabel metal2 s 139660 158648 139716 159448 6 m_in[227]
port 143 nsew signal input
rlabel metal2 s 140212 158648 140268 159448 6 m_in[228]
port 144 nsew signal input
rlabel metal2 s 140856 158648 140912 159448 6 m_in[229]
port 145 nsew signal input
rlabel metal2 s 13528 158648 13584 159448 6 m_in[22]
port 146 nsew signal input
rlabel metal2 s 141500 158648 141556 159448 6 m_in[230]
port 147 nsew signal input
rlabel metal2 s 142144 158648 142200 159448 6 m_in[231]
port 148 nsew signal input
rlabel metal2 s 142696 158648 142752 159448 6 m_in[232]
port 149 nsew signal input
rlabel metal2 s 143340 158648 143396 159448 6 m_in[233]
port 150 nsew signal input
rlabel metal2 s 143984 158648 144040 159448 6 m_in[234]
port 151 nsew signal input
rlabel metal2 s 144536 158648 144592 159448 6 m_in[235]
port 152 nsew signal input
rlabel metal2 s 145180 158648 145236 159448 6 m_in[236]
port 153 nsew signal input
rlabel metal2 s 145824 158648 145880 159448 6 m_in[237]
port 154 nsew signal input
rlabel metal2 s 146376 158648 146432 159448 6 m_in[238]
port 155 nsew signal input
rlabel metal2 s 147020 158648 147076 159448 6 m_in[239]
port 156 nsew signal input
rlabel metal2 s 14080 158648 14136 159448 6 m_in[23]
port 157 nsew signal input
rlabel metal2 s 147664 158648 147720 159448 6 m_in[240]
port 158 nsew signal input
rlabel metal2 s 148216 158648 148272 159448 6 m_in[241]
port 159 nsew signal input
rlabel metal2 s 148860 158648 148916 159448 6 m_in[242]
port 160 nsew signal input
rlabel metal2 s 149504 158648 149560 159448 6 m_in[243]
port 161 nsew signal input
rlabel metal2 s 150056 158648 150112 159448 6 m_in[244]
port 162 nsew signal input
rlabel metal2 s 150700 158648 150756 159448 6 m_in[245]
port 163 nsew signal input
rlabel metal2 s 151344 158648 151400 159448 6 m_in[246]
port 164 nsew signal input
rlabel metal2 s 151988 158648 152044 159448 6 m_in[247]
port 165 nsew signal input
rlabel metal2 s 152540 158648 152596 159448 6 m_in[248]
port 166 nsew signal input
rlabel metal2 s 153184 158648 153240 159448 6 m_in[249]
port 167 nsew signal input
rlabel metal2 s 14724 158648 14780 159448 6 m_in[24]
port 168 nsew signal input
rlabel metal2 s 153828 158648 153884 159448 6 m_in[250]
port 169 nsew signal input
rlabel metal2 s 154380 158648 154436 159448 6 m_in[251]
port 170 nsew signal input
rlabel metal2 s 155024 158648 155080 159448 6 m_in[252]
port 171 nsew signal input
rlabel metal2 s 155668 158648 155724 159448 6 m_in[253]
port 172 nsew signal input
rlabel metal2 s 156220 158648 156276 159448 6 m_in[254]
port 173 nsew signal input
rlabel metal2 s 156864 158648 156920 159448 6 m_in[255]
port 174 nsew signal input
rlabel metal2 s 157508 158648 157564 159448 6 m_in[256]
port 175 nsew signal input
rlabel metal2 s 158060 158648 158116 159448 6 m_in[257]
port 176 nsew signal input
rlabel metal2 s 158704 158648 158760 159448 6 m_in[258]
port 177 nsew signal input
rlabel metal2 s 15368 158648 15424 159448 6 m_in[25]
port 178 nsew signal input
rlabel metal2 s 15920 158648 15976 159448 6 m_in[26]
port 179 nsew signal input
rlabel metal2 s 16564 158648 16620 159448 6 m_in[27]
port 180 nsew signal input
rlabel metal2 s 17208 158648 17264 159448 6 m_in[28]
port 181 nsew signal input
rlabel metal2 s 17760 158648 17816 159448 6 m_in[29]
port 182 nsew signal input
rlabel metal2 s 1200 158648 1256 159448 6 m_in[2]
port 183 nsew signal input
rlabel metal2 s 18404 158648 18460 159448 6 m_in[30]
port 184 nsew signal input
rlabel metal2 s 19048 158648 19104 159448 6 m_in[31]
port 185 nsew signal input
rlabel metal2 s 19692 158648 19748 159448 6 m_in[32]
port 186 nsew signal input
rlabel metal2 s 20244 158648 20300 159448 6 m_in[33]
port 187 nsew signal input
rlabel metal2 s 20888 158648 20944 159448 6 m_in[34]
port 188 nsew signal input
rlabel metal2 s 21532 158648 21588 159448 6 m_in[35]
port 189 nsew signal input
rlabel metal2 s 22084 158648 22140 159448 6 m_in[36]
port 190 nsew signal input
rlabel metal2 s 22728 158648 22784 159448 6 m_in[37]
port 191 nsew signal input
rlabel metal2 s 23372 158648 23428 159448 6 m_in[38]
port 192 nsew signal input
rlabel metal2 s 23924 158648 23980 159448 6 m_in[39]
port 193 nsew signal input
rlabel metal2 s 1844 158648 1900 159448 6 m_in[3]
port 194 nsew signal input
rlabel metal2 s 24568 158648 24624 159448 6 m_in[40]
port 195 nsew signal input
rlabel metal2 s 25212 158648 25268 159448 6 m_in[41]
port 196 nsew signal input
rlabel metal2 s 25764 158648 25820 159448 6 m_in[42]
port 197 nsew signal input
rlabel metal2 s 26408 158648 26464 159448 6 m_in[43]
port 198 nsew signal input
rlabel metal2 s 27052 158648 27108 159448 6 m_in[44]
port 199 nsew signal input
rlabel metal2 s 27604 158648 27660 159448 6 m_in[45]
port 200 nsew signal input
rlabel metal2 s 28248 158648 28304 159448 6 m_in[46]
port 201 nsew signal input
rlabel metal2 s 28892 158648 28948 159448 6 m_in[47]
port 202 nsew signal input
rlabel metal2 s 29536 158648 29592 159448 6 m_in[48]
port 203 nsew signal input
rlabel metal2 s 30088 158648 30144 159448 6 m_in[49]
port 204 nsew signal input
rlabel metal2 s 2396 158648 2452 159448 6 m_in[4]
port 205 nsew signal input
rlabel metal2 s 30732 158648 30788 159448 6 m_in[50]
port 206 nsew signal input
rlabel metal2 s 31376 158648 31432 159448 6 m_in[51]
port 207 nsew signal input
rlabel metal2 s 31928 158648 31984 159448 6 m_in[52]
port 208 nsew signal input
rlabel metal2 s 32572 158648 32628 159448 6 m_in[53]
port 209 nsew signal input
rlabel metal2 s 33216 158648 33272 159448 6 m_in[54]
port 210 nsew signal input
rlabel metal2 s 33768 158648 33824 159448 6 m_in[55]
port 211 nsew signal input
rlabel metal2 s 34412 158648 34468 159448 6 m_in[56]
port 212 nsew signal input
rlabel metal2 s 35056 158648 35112 159448 6 m_in[57]
port 213 nsew signal input
rlabel metal2 s 35608 158648 35664 159448 6 m_in[58]
port 214 nsew signal input
rlabel metal2 s 36252 158648 36308 159448 6 m_in[59]
port 215 nsew signal input
rlabel metal2 s 3040 158648 3096 159448 6 m_in[5]
port 216 nsew signal input
rlabel metal2 s 36896 158648 36952 159448 6 m_in[60]
port 217 nsew signal input
rlabel metal2 s 37448 158648 37504 159448 6 m_in[61]
port 218 nsew signal input
rlabel metal2 s 38092 158648 38148 159448 6 m_in[62]
port 219 nsew signal input
rlabel metal2 s 38736 158648 38792 159448 6 m_in[63]
port 220 nsew signal input
rlabel metal2 s 39380 158648 39436 159448 6 m_in[64]
port 221 nsew signal input
rlabel metal2 s 39932 158648 39988 159448 6 m_in[65]
port 222 nsew signal input
rlabel metal2 s 40576 158648 40632 159448 6 m_in[66]
port 223 nsew signal input
rlabel metal2 s 41220 158648 41276 159448 6 m_in[67]
port 224 nsew signal input
rlabel metal2 s 41772 158648 41828 159448 6 m_in[68]
port 225 nsew signal input
rlabel metal2 s 42416 158648 42472 159448 6 m_in[69]
port 226 nsew signal input
rlabel metal2 s 3684 158648 3740 159448 6 m_in[6]
port 227 nsew signal input
rlabel metal2 s 43060 158648 43116 159448 6 m_in[70]
port 228 nsew signal input
rlabel metal2 s 43612 158648 43668 159448 6 m_in[71]
port 229 nsew signal input
rlabel metal2 s 44256 158648 44312 159448 6 m_in[72]
port 230 nsew signal input
rlabel metal2 s 44900 158648 44956 159448 6 m_in[73]
port 231 nsew signal input
rlabel metal2 s 45452 158648 45508 159448 6 m_in[74]
port 232 nsew signal input
rlabel metal2 s 46096 158648 46152 159448 6 m_in[75]
port 233 nsew signal input
rlabel metal2 s 46740 158648 46796 159448 6 m_in[76]
port 234 nsew signal input
rlabel metal2 s 47384 158648 47440 159448 6 m_in[77]
port 235 nsew signal input
rlabel metal2 s 47936 158648 47992 159448 6 m_in[78]
port 236 nsew signal input
rlabel metal2 s 48580 158648 48636 159448 6 m_in[79]
port 237 nsew signal input
rlabel metal2 s 4236 158648 4292 159448 6 m_in[7]
port 238 nsew signal input
rlabel metal2 s 49224 158648 49280 159448 6 m_in[80]
port 239 nsew signal input
rlabel metal2 s 49776 158648 49832 159448 6 m_in[81]
port 240 nsew signal input
rlabel metal2 s 50420 158648 50476 159448 6 m_in[82]
port 241 nsew signal input
rlabel metal2 s 51064 158648 51120 159448 6 m_in[83]
port 242 nsew signal input
rlabel metal2 s 51616 158648 51672 159448 6 m_in[84]
port 243 nsew signal input
rlabel metal2 s 52260 158648 52316 159448 6 m_in[85]
port 244 nsew signal input
rlabel metal2 s 52904 158648 52960 159448 6 m_in[86]
port 245 nsew signal input
rlabel metal2 s 53456 158648 53512 159448 6 m_in[87]
port 246 nsew signal input
rlabel metal2 s 54100 158648 54156 159448 6 m_in[88]
port 247 nsew signal input
rlabel metal2 s 54744 158648 54800 159448 6 m_in[89]
port 248 nsew signal input
rlabel metal2 s 4880 158648 4936 159448 6 m_in[8]
port 249 nsew signal input
rlabel metal2 s 55296 158648 55352 159448 6 m_in[90]
port 250 nsew signal input
rlabel metal2 s 55940 158648 55996 159448 6 m_in[91]
port 251 nsew signal input
rlabel metal2 s 56584 158648 56640 159448 6 m_in[92]
port 252 nsew signal input
rlabel metal2 s 57228 158648 57284 159448 6 m_in[93]
port 253 nsew signal input
rlabel metal2 s 57780 158648 57836 159448 6 m_in[94]
port 254 nsew signal input
rlabel metal2 s 58424 158648 58480 159448 6 m_in[95]
port 255 nsew signal input
rlabel metal2 s 59068 158648 59124 159448 6 m_in[96]
port 256 nsew signal input
rlabel metal2 s 59620 158648 59676 159448 6 m_in[97]
port 257 nsew signal input
rlabel metal2 s 60264 158648 60320 159448 6 m_in[98]
port 258 nsew signal input
rlabel metal2 s 60908 158648 60964 159448 6 m_in[99]
port 259 nsew signal input
rlabel metal2 s 5524 158648 5580 159448 6 m_in[9]
port 260 nsew signal input
rlabel metal3 s 158910 0 159710 120 6 m_out[0]
port 261 nsew signal output
rlabel metal3 s 158910 122944 159710 123064 6 m_out[100]
port 262 nsew signal output
rlabel metal3 s 158910 124168 159710 124288 6 m_out[101]
port 263 nsew signal output
rlabel metal3 s 158910 125392 159710 125512 6 m_out[102]
port 264 nsew signal output
rlabel metal3 s 158910 126616 159710 126736 6 m_out[103]
port 265 nsew signal output
rlabel metal3 s 158910 127840 159710 127960 6 m_out[104]
port 266 nsew signal output
rlabel metal3 s 158910 129064 159710 129184 6 m_out[105]
port 267 nsew signal output
rlabel metal3 s 158910 130288 159710 130408 6 m_out[106]
port 268 nsew signal output
rlabel metal3 s 158910 131512 159710 131632 6 m_out[107]
port 269 nsew signal output
rlabel metal3 s 158910 132736 159710 132856 6 m_out[108]
port 270 nsew signal output
rlabel metal3 s 158910 134096 159710 134216 6 m_out[109]
port 271 nsew signal output
rlabel metal3 s 158910 12240 159710 12360 6 m_out[10]
port 272 nsew signal output
rlabel metal3 s 158910 135320 159710 135440 6 m_out[110]
port 273 nsew signal output
rlabel metal3 s 158910 136544 159710 136664 6 m_out[111]
port 274 nsew signal output
rlabel metal3 s 158910 137768 159710 137888 6 m_out[112]
port 275 nsew signal output
rlabel metal3 s 158910 138992 159710 139112 6 m_out[113]
port 276 nsew signal output
rlabel metal3 s 158910 140216 159710 140336 6 m_out[114]
port 277 nsew signal output
rlabel metal3 s 158910 141440 159710 141560 6 m_out[115]
port 278 nsew signal output
rlabel metal3 s 158910 142664 159710 142784 6 m_out[116]
port 279 nsew signal output
rlabel metal3 s 158910 143888 159710 144008 6 m_out[117]
port 280 nsew signal output
rlabel metal3 s 158910 145112 159710 145232 6 m_out[118]
port 281 nsew signal output
rlabel metal3 s 158910 146336 159710 146456 6 m_out[119]
port 282 nsew signal output
rlabel metal3 s 158910 13464 159710 13584 6 m_out[11]
port 283 nsew signal output
rlabel metal3 s 158910 147560 159710 147680 6 m_out[120]
port 284 nsew signal output
rlabel metal3 s 158910 148784 159710 148904 6 m_out[121]
port 285 nsew signal output
rlabel metal3 s 158910 150008 159710 150128 6 m_out[122]
port 286 nsew signal output
rlabel metal3 s 158910 151232 159710 151352 6 m_out[123]
port 287 nsew signal output
rlabel metal3 s 158910 152456 159710 152576 6 m_out[124]
port 288 nsew signal output
rlabel metal3 s 158910 153680 159710 153800 6 m_out[125]
port 289 nsew signal output
rlabel metal3 s 158910 154904 159710 155024 6 m_out[126]
port 290 nsew signal output
rlabel metal3 s 158910 156128 159710 156248 6 m_out[127]
port 291 nsew signal output
rlabel metal3 s 158910 157352 159710 157472 6 m_out[128]
port 292 nsew signal output
rlabel metal3 s 158910 158576 159710 158696 6 m_out[129]
port 293 nsew signal output
rlabel metal3 s 158910 14688 159710 14808 6 m_out[12]
port 294 nsew signal output
rlabel metal3 s 158910 15912 159710 16032 6 m_out[13]
port 295 nsew signal output
rlabel metal3 s 158910 17136 159710 17256 6 m_out[14]
port 296 nsew signal output
rlabel metal3 s 158910 18360 159710 18480 6 m_out[15]
port 297 nsew signal output
rlabel metal3 s 158910 19584 159710 19704 6 m_out[16]
port 298 nsew signal output
rlabel metal3 s 158910 20808 159710 20928 6 m_out[17]
port 299 nsew signal output
rlabel metal3 s 158910 22032 159710 22152 6 m_out[18]
port 300 nsew signal output
rlabel metal3 s 158910 23256 159710 23376 6 m_out[19]
port 301 nsew signal output
rlabel metal3 s 158910 1224 159710 1344 6 m_out[1]
port 302 nsew signal output
rlabel metal3 s 158910 24480 159710 24600 6 m_out[20]
port 303 nsew signal output
rlabel metal3 s 158910 25704 159710 25824 6 m_out[21]
port 304 nsew signal output
rlabel metal3 s 158910 27064 159710 27184 6 m_out[22]
port 305 nsew signal output
rlabel metal3 s 158910 28288 159710 28408 6 m_out[23]
port 306 nsew signal output
rlabel metal3 s 158910 29512 159710 29632 6 m_out[24]
port 307 nsew signal output
rlabel metal3 s 158910 30736 159710 30856 6 m_out[25]
port 308 nsew signal output
rlabel metal3 s 158910 31960 159710 32080 6 m_out[26]
port 309 nsew signal output
rlabel metal3 s 158910 33184 159710 33304 6 m_out[27]
port 310 nsew signal output
rlabel metal3 s 158910 34408 159710 34528 6 m_out[28]
port 311 nsew signal output
rlabel metal3 s 158910 35632 159710 35752 6 m_out[29]
port 312 nsew signal output
rlabel metal3 s 158910 2448 159710 2568 6 m_out[2]
port 313 nsew signal output
rlabel metal3 s 158910 36856 159710 36976 6 m_out[30]
port 314 nsew signal output
rlabel metal3 s 158910 38080 159710 38200 6 m_out[31]
port 315 nsew signal output
rlabel metal3 s 158910 39304 159710 39424 6 m_out[32]
port 316 nsew signal output
rlabel metal3 s 158910 40528 159710 40648 6 m_out[33]
port 317 nsew signal output
rlabel metal3 s 158910 41752 159710 41872 6 m_out[34]
port 318 nsew signal output
rlabel metal3 s 158910 42976 159710 43096 6 m_out[35]
port 319 nsew signal output
rlabel metal3 s 158910 44200 159710 44320 6 m_out[36]
port 320 nsew signal output
rlabel metal3 s 158910 45424 159710 45544 6 m_out[37]
port 321 nsew signal output
rlabel metal3 s 158910 46648 159710 46768 6 m_out[38]
port 322 nsew signal output
rlabel metal3 s 158910 47872 159710 47992 6 m_out[39]
port 323 nsew signal output
rlabel metal3 s 158910 3672 159710 3792 6 m_out[3]
port 324 nsew signal output
rlabel metal3 s 158910 49096 159710 49216 6 m_out[40]
port 325 nsew signal output
rlabel metal3 s 158910 50320 159710 50440 6 m_out[41]
port 326 nsew signal output
rlabel metal3 s 158910 51544 159710 51664 6 m_out[42]
port 327 nsew signal output
rlabel metal3 s 158910 52768 159710 52888 6 m_out[43]
port 328 nsew signal output
rlabel metal3 s 158910 54128 159710 54248 6 m_out[44]
port 329 nsew signal output
rlabel metal3 s 158910 55352 159710 55472 6 m_out[45]
port 330 nsew signal output
rlabel metal3 s 158910 56576 159710 56696 6 m_out[46]
port 331 nsew signal output
rlabel metal3 s 158910 57800 159710 57920 6 m_out[47]
port 332 nsew signal output
rlabel metal3 s 158910 59024 159710 59144 6 m_out[48]
port 333 nsew signal output
rlabel metal3 s 158910 60248 159710 60368 6 m_out[49]
port 334 nsew signal output
rlabel metal3 s 158910 4896 159710 5016 6 m_out[4]
port 335 nsew signal output
rlabel metal3 s 158910 61472 159710 61592 6 m_out[50]
port 336 nsew signal output
rlabel metal3 s 158910 62696 159710 62816 6 m_out[51]
port 337 nsew signal output
rlabel metal3 s 158910 63920 159710 64040 6 m_out[52]
port 338 nsew signal output
rlabel metal3 s 158910 65144 159710 65264 6 m_out[53]
port 339 nsew signal output
rlabel metal3 s 158910 66368 159710 66488 6 m_out[54]
port 340 nsew signal output
rlabel metal3 s 158910 67592 159710 67712 6 m_out[55]
port 341 nsew signal output
rlabel metal3 s 158910 68816 159710 68936 6 m_out[56]
port 342 nsew signal output
rlabel metal3 s 158910 70040 159710 70160 6 m_out[57]
port 343 nsew signal output
rlabel metal3 s 158910 71264 159710 71384 6 m_out[58]
port 344 nsew signal output
rlabel metal3 s 158910 72488 159710 72608 6 m_out[59]
port 345 nsew signal output
rlabel metal3 s 158910 6120 159710 6240 6 m_out[5]
port 346 nsew signal output
rlabel metal3 s 158910 73712 159710 73832 6 m_out[60]
port 347 nsew signal output
rlabel metal3 s 158910 74936 159710 75056 6 m_out[61]
port 348 nsew signal output
rlabel metal3 s 158910 76160 159710 76280 6 m_out[62]
port 349 nsew signal output
rlabel metal3 s 158910 77384 159710 77504 6 m_out[63]
port 350 nsew signal output
rlabel metal3 s 158910 78608 159710 78728 6 m_out[64]
port 351 nsew signal output
rlabel metal3 s 158910 79968 159710 80088 6 m_out[65]
port 352 nsew signal output
rlabel metal3 s 158910 81192 159710 81312 6 m_out[66]
port 353 nsew signal output
rlabel metal3 s 158910 82416 159710 82536 6 m_out[67]
port 354 nsew signal output
rlabel metal3 s 158910 83640 159710 83760 6 m_out[68]
port 355 nsew signal output
rlabel metal3 s 158910 84864 159710 84984 6 m_out[69]
port 356 nsew signal output
rlabel metal3 s 158910 7344 159710 7464 6 m_out[6]
port 357 nsew signal output
rlabel metal3 s 158910 86088 159710 86208 6 m_out[70]
port 358 nsew signal output
rlabel metal3 s 158910 87312 159710 87432 6 m_out[71]
port 359 nsew signal output
rlabel metal3 s 158910 88536 159710 88656 6 m_out[72]
port 360 nsew signal output
rlabel metal3 s 158910 89760 159710 89880 6 m_out[73]
port 361 nsew signal output
rlabel metal3 s 158910 90984 159710 91104 6 m_out[74]
port 362 nsew signal output
rlabel metal3 s 158910 92208 159710 92328 6 m_out[75]
port 363 nsew signal output
rlabel metal3 s 158910 93432 159710 93552 6 m_out[76]
port 364 nsew signal output
rlabel metal3 s 158910 94656 159710 94776 6 m_out[77]
port 365 nsew signal output
rlabel metal3 s 158910 95880 159710 96000 6 m_out[78]
port 366 nsew signal output
rlabel metal3 s 158910 97104 159710 97224 6 m_out[79]
port 367 nsew signal output
rlabel metal3 s 158910 8568 159710 8688 6 m_out[7]
port 368 nsew signal output
rlabel metal3 s 158910 98328 159710 98448 6 m_out[80]
port 369 nsew signal output
rlabel metal3 s 158910 99552 159710 99672 6 m_out[81]
port 370 nsew signal output
rlabel metal3 s 158910 100776 159710 100896 6 m_out[82]
port 371 nsew signal output
rlabel metal3 s 158910 102000 159710 102120 6 m_out[83]
port 372 nsew signal output
rlabel metal3 s 158910 103224 159710 103344 6 m_out[84]
port 373 nsew signal output
rlabel metal3 s 158910 104448 159710 104568 6 m_out[85]
port 374 nsew signal output
rlabel metal3 s 158910 105672 159710 105792 6 m_out[86]
port 375 nsew signal output
rlabel metal3 s 158910 107032 159710 107152 6 m_out[87]
port 376 nsew signal output
rlabel metal3 s 158910 108256 159710 108376 6 m_out[88]
port 377 nsew signal output
rlabel metal3 s 158910 109480 159710 109600 6 m_out[89]
port 378 nsew signal output
rlabel metal3 s 158910 9792 159710 9912 6 m_out[8]
port 379 nsew signal output
rlabel metal3 s 158910 110704 159710 110824 6 m_out[90]
port 380 nsew signal output
rlabel metal3 s 158910 111928 159710 112048 6 m_out[91]
port 381 nsew signal output
rlabel metal3 s 158910 113152 159710 113272 6 m_out[92]
port 382 nsew signal output
rlabel metal3 s 158910 114376 159710 114496 6 m_out[93]
port 383 nsew signal output
rlabel metal3 s 158910 115600 159710 115720 6 m_out[94]
port 384 nsew signal output
rlabel metal3 s 158910 116824 159710 116944 6 m_out[95]
port 385 nsew signal output
rlabel metal3 s 158910 118048 159710 118168 6 m_out[96]
port 386 nsew signal output
rlabel metal3 s 158910 119272 159710 119392 6 m_out[97]
port 387 nsew signal output
rlabel metal3 s 158910 120496 159710 120616 6 m_out[98]
port 388 nsew signal output
rlabel metal3 s 158910 121720 159710 121840 6 m_out[99]
port 389 nsew signal output
rlabel metal3 s 158910 11016 159710 11136 6 m_out[9]
port 390 nsew signal output
rlabel metal4 s 157518 1576 157838 157256 6 vccd1
port 391 nsew power bidirectional
rlabel metal4 s 126798 1576 127118 157256 6 vccd1
port 392 nsew power bidirectional
rlabel metal4 s 96078 1576 96398 157256 6 vccd1
port 393 nsew power bidirectional
rlabel metal4 s 65358 1576 65678 157256 6 vccd1
port 394 nsew power bidirectional
rlabel metal4 s 34638 1576 34958 157256 6 vccd1
port 395 nsew power bidirectional
rlabel metal4 s 3918 1576 4238 157256 6 vccd1
port 396 nsew power bidirectional
rlabel metal4 s 142158 1576 142478 157256 6 vssd1
port 397 nsew ground bidirectional
rlabel metal4 s 111438 1576 111758 157256 6 vssd1
port 398 nsew ground bidirectional
rlabel metal4 s 80718 1576 81038 157256 6 vssd1
port 399 nsew ground bidirectional
rlabel metal4 s 49998 1576 50318 157256 6 vssd1
port 400 nsew ground bidirectional
rlabel metal4 s 19278 1576 19598 157256 6 vssd1
port 401 nsew ground bidirectional
rlabel metal4 s 127458 1624 127778 157208 6 vccd2
port 402 nsew power bidirectional
rlabel metal4 s 96738 1624 97058 157208 6 vccd2
port 403 nsew power bidirectional
rlabel metal4 s 66018 1624 66338 157208 6 vccd2
port 404 nsew power bidirectional
rlabel metal4 s 35298 1624 35618 157208 6 vccd2
port 405 nsew power bidirectional
rlabel metal4 s 4578 1624 4898 157208 6 vccd2
port 406 nsew power bidirectional
rlabel metal4 s 142818 1624 143138 157208 6 vssd2
port 407 nsew ground bidirectional
rlabel metal4 s 112098 1624 112418 157208 6 vssd2
port 408 nsew ground bidirectional
rlabel metal4 s 81378 1624 81698 157208 6 vssd2
port 409 nsew ground bidirectional
rlabel metal4 s 50658 1624 50978 157208 6 vssd2
port 410 nsew ground bidirectional
rlabel metal4 s 19938 1624 20258 157208 6 vssd2
port 411 nsew ground bidirectional
rlabel metal4 s 128118 1624 128438 157208 6 vdda1
port 412 nsew power bidirectional
rlabel metal4 s 97398 1624 97718 157208 6 vdda1
port 413 nsew power bidirectional
rlabel metal4 s 66678 1624 66998 157208 6 vdda1
port 414 nsew power bidirectional
rlabel metal4 s 35958 1624 36278 157208 6 vdda1
port 415 nsew power bidirectional
rlabel metal4 s 5238 1624 5558 157208 6 vdda1
port 416 nsew power bidirectional
rlabel metal4 s 143478 1624 143798 157208 6 vssa1
port 417 nsew ground bidirectional
rlabel metal4 s 112758 1624 113078 157208 6 vssa1
port 418 nsew ground bidirectional
rlabel metal4 s 82038 1624 82358 157208 6 vssa1
port 419 nsew ground bidirectional
rlabel metal4 s 51318 1624 51638 157208 6 vssa1
port 420 nsew ground bidirectional
rlabel metal4 s 20598 1624 20918 157208 6 vssa1
port 421 nsew ground bidirectional
rlabel metal4 s 128778 1624 129098 157208 6 vdda2
port 422 nsew power bidirectional
rlabel metal4 s 98058 1624 98378 157208 6 vdda2
port 423 nsew power bidirectional
rlabel metal4 s 67338 1624 67658 157208 6 vdda2
port 424 nsew power bidirectional
rlabel metal4 s 36618 1624 36938 157208 6 vdda2
port 425 nsew power bidirectional
rlabel metal4 s 5898 1624 6218 157208 6 vdda2
port 426 nsew power bidirectional
rlabel metal4 s 144138 1624 144458 157208 6 vssa2
port 427 nsew ground bidirectional
rlabel metal4 s 113418 1624 113738 157208 6 vssa2
port 428 nsew ground bidirectional
rlabel metal4 s 82698 1624 83018 157208 6 vssa2
port 429 nsew ground bidirectional
rlabel metal4 s 51978 1624 52298 157208 6 vssa2
port 430 nsew ground bidirectional
rlabel metal4 s 21258 1624 21578 157208 6 vssa2
port 431 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 159710 159448
string LEFview TRUE
<< end >>
