magic
tech sky130A
magscale 1 2
timestamp 1610963659
<< nwell >>
rect 0 117231 577836 117542
rect 0 117221 206317 117231
rect 0 116689 74757 116699
rect 0 116143 577836 116689
rect 0 116133 62245 116143
rect 0 115601 12841 115611
rect 0 115055 577836 115601
rect 0 115045 7689 115055
rect 0 114513 25629 114523
rect 0 113967 577836 114513
rect 0 113957 14773 113967
rect 0 113425 24249 113435
rect 0 112879 577836 113425
rect 0 112869 15785 112879
rect 0 112337 15049 112347
rect 0 111791 577836 112337
rect 0 111781 4193 111791
rect 0 111249 3641 111259
rect 0 110703 577836 111249
rect 0 110693 21397 110703
rect 0 110161 16521 110171
rect 0 109615 577836 110161
rect 0 109605 52769 109615
rect 0 109073 23513 109083
rect 0 108527 577836 109073
rect 0 108517 11553 108527
rect 0 107985 55161 107995
rect 0 107439 577836 107985
rect 0 107429 4377 107439
rect 0 106897 8793 106907
rect 0 106351 577836 106897
rect 0 106341 50837 106351
rect 0 105809 13025 105819
rect 0 105263 577836 105809
rect 0 105253 12565 105263
rect 0 104721 8793 104731
rect 0 104175 577836 104721
rect 0 104165 35749 104175
rect 0 103633 14497 103643
rect 0 103087 577836 103633
rect 0 103077 21397 103087
rect 0 102545 7137 102555
rect 0 101999 577836 102545
rect 0 101989 18637 101999
rect 0 101457 10541 101467
rect 0 100911 577836 101457
rect 0 100901 6493 100911
rect 0 100369 79449 100379
rect 0 99823 577836 100369
rect 0 99813 4193 99823
rect 0 99281 3181 99291
rect 0 98735 577836 99281
rect 0 98725 42649 98735
rect 0 98193 59301 98203
rect 0 97647 577836 98193
rect 0 97637 11553 97647
rect 0 97105 6401 97115
rect 0 96559 577836 97105
rect 0 96549 49457 96559
rect 0 96017 7321 96027
rect 0 95471 577836 96017
rect 0 95461 42097 95471
rect 0 94929 16245 94939
rect 0 94383 577836 94929
rect 0 94373 25169 94383
rect 0 93841 15601 93851
rect 0 93295 577836 93841
rect 0 93285 17165 93295
rect 0 92753 5389 92763
rect 0 92207 577836 92753
rect 0 92197 41821 92207
rect 0 91665 12565 91675
rect 0 91119 577836 91665
rect 0 91109 3365 91119
rect 0 90577 3181 90587
rect 0 90031 577836 90577
rect 0 90021 84509 90031
rect 0 89489 37221 89499
rect 0 88943 577836 89489
rect 0 88933 42097 88943
rect 0 88401 7045 88411
rect 0 87855 577836 88401
rect 0 87845 11553 87855
rect 0 87313 18637 87323
rect 0 86767 577836 87313
rect 0 86757 45225 86767
rect 0 86225 31885 86235
rect 0 85679 577836 86225
rect 0 85669 39797 85679
rect 0 85137 18637 85147
rect 0 84591 577836 85137
rect 0 84581 49089 84591
rect 0 84049 7229 84059
rect 0 83503 577836 84049
rect 0 83493 29125 83503
rect 0 82961 11553 82971
rect 0 82415 577836 82961
rect 0 82405 9713 82415
rect 0 81873 39061 81883
rect 0 81327 577836 81873
rect 0 81317 9529 81327
rect 0 80785 28481 80795
rect 0 80239 577836 80785
rect 0 80229 17165 80239
rect 0 79697 38049 79707
rect 0 79151 577836 79697
rect 0 79141 17165 79151
rect 0 78609 14405 78619
rect 0 78063 577836 78609
rect 0 78053 68593 78063
rect 0 77521 3181 77531
rect 0 76975 577836 77521
rect 0 76965 22777 76975
rect 0 76433 6033 76443
rect 0 75887 577836 76433
rect 0 75877 67673 75887
rect 0 75345 13025 75355
rect 0 74799 577836 75345
rect 0 74789 52861 74799
rect 0 74257 8793 74267
rect 0 73711 577836 74257
rect 0 73701 17165 73711
rect 0 73169 6861 73179
rect 0 72623 577836 73169
rect 0 72613 28389 72623
rect 0 72081 3181 72091
rect 0 71535 577836 72081
rect 0 71525 30689 71535
rect 0 70993 513 71003
rect 0 70447 577836 70993
rect 0 70437 131061 70447
rect 0 69905 3181 69915
rect 0 69359 577836 69905
rect 0 69349 3273 69359
rect 0 68817 14865 68827
rect 0 68271 577836 68817
rect 0 68261 15233 68271
rect 0 67729 22317 67739
rect 0 67183 577836 67729
rect 0 67173 1157 67183
rect 0 66641 7229 66651
rect 0 66095 577836 66641
rect 0 66085 1525 66095
rect 0 65553 3181 65563
rect 0 65007 577836 65553
rect 0 64997 45317 65007
rect 0 64465 20017 64475
rect 0 63919 577836 64465
rect 0 63909 19281 63919
rect 0 63377 36853 63387
rect 0 62831 577836 63377
rect 0 62821 2537 62831
rect 0 62289 46513 62299
rect 0 61743 577836 62289
rect 0 61733 1341 61743
rect 0 61201 46697 61211
rect 0 60655 577836 61201
rect 0 60645 25445 60655
rect 0 60113 1525 60123
rect 0 59567 577836 60113
rect 0 59557 34001 59567
rect 0 59025 42465 59035
rect 0 58479 577836 59025
rect 0 58469 51297 58479
rect 0 57937 110545 57947
rect 0 57391 577836 57937
rect 0 57381 2629 57391
rect 0 56849 9345 56859
rect 0 56303 577836 56849
rect 0 56293 48353 56303
rect 0 55761 29217 55771
rect 0 55215 577836 55761
rect 0 55205 2537 55215
rect 0 54673 60773 54683
rect 0 54127 577836 54673
rect 0 54117 15785 54127
rect 0 53585 6401 53595
rect 0 53039 577836 53585
rect 0 53029 3641 53039
rect 0 52497 12105 52507
rect 0 51951 577836 52497
rect 0 51941 37313 51951
rect 0 51409 28665 51419
rect 0 50863 577836 51409
rect 0 50853 13393 50863
rect 0 50321 15877 50331
rect 0 49775 577836 50321
rect 0 49765 1157 49775
rect 0 49233 84785 49243
rect 0 48687 577836 49233
rect 0 48677 14589 48687
rect 0 48145 12933 48155
rect 0 47599 577836 48145
rect 0 47589 11553 47599
rect 0 47057 5113 47067
rect 0 46511 577836 47057
rect 0 46501 59853 46511
rect 0 45969 17993 45979
rect 0 45423 577836 45969
rect 0 45413 6861 45423
rect 0 44881 121953 44891
rect 0 44335 577836 44881
rect 0 44325 83129 44335
rect 0 43793 39061 43803
rect 0 43247 577836 43793
rect 0 43237 24893 43247
rect 0 42705 10081 42715
rect 0 42159 577836 42705
rect 0 42149 24341 42159
rect 0 41617 40441 41627
rect 0 41071 577836 41617
rect 0 41061 3365 41071
rect 0 40529 27745 40539
rect 0 39983 577836 40529
rect 0 39973 3549 39983
rect 0 39441 10817 39451
rect 0 38895 577836 39441
rect 0 38885 25261 38895
rect 0 38353 20017 38363
rect 0 37807 577836 38353
rect 0 37797 17165 37807
rect 0 37265 37865 37275
rect 0 36719 577836 37265
rect 0 36709 23789 36719
rect 0 36177 38601 36187
rect 0 35631 577836 36177
rect 0 35621 605 35631
rect 0 35089 4193 35099
rect 0 34543 577836 35089
rect 0 34533 13025 34543
rect 0 34001 8793 34011
rect 0 33455 577836 34001
rect 0 33445 1617 33455
rect 0 32913 1801 32923
rect 0 32367 577836 32913
rect 0 32357 5941 32367
rect 0 31825 48077 31835
rect 0 31279 577836 31825
rect 0 31269 47709 31279
rect 0 30737 70525 30747
rect 0 30191 577836 30737
rect 0 30181 224809 30191
rect 0 29649 10817 29659
rect 0 29103 577836 29649
rect 0 29093 6309 29103
rect 0 28561 6125 28571
rect 0 28015 577836 28561
rect 0 28005 18637 28015
rect 0 27473 32805 27483
rect 0 26927 577836 27473
rect 0 26917 11553 26927
rect 0 26385 36853 26395
rect 0 25839 577836 26385
rect 0 25829 34737 25839
rect 0 25297 11277 25307
rect 0 24751 577836 25297
rect 0 24741 87913 24751
rect 0 24209 11093 24219
rect 0 23663 577836 24209
rect 0 23653 11553 23663
rect 0 23121 35473 23131
rect 0 22575 577836 23121
rect 0 22565 13669 22575
rect 0 22033 44489 22043
rect 0 21487 577836 22033
rect 0 21477 9713 21487
rect 0 20945 6585 20955
rect 0 20399 577836 20945
rect 0 20389 34553 20399
rect 0 19857 7321 19867
rect 0 19311 577836 19857
rect 0 19301 15693 19311
rect 0 18769 151761 18779
rect 0 18223 577836 18769
rect 0 18213 2997 18223
rect 0 17681 35289 17691
rect 0 17135 577836 17681
rect 0 17125 37405 17135
rect 0 16593 16889 16603
rect 0 16047 577836 16593
rect 0 16037 52861 16047
rect 0 15505 22777 15515
rect 0 14959 577836 15505
rect 0 14949 24157 14959
rect 0 14417 11185 14427
rect 0 13871 577836 14417
rect 0 13861 28849 13871
rect 0 13329 3365 13339
rect 0 12783 577836 13329
rect 0 12773 47525 12783
rect 0 12241 44029 12251
rect 0 11695 577836 12241
rect 0 11685 11553 11695
rect 0 11153 10817 11163
rect 0 10607 577836 11153
rect 0 10597 68409 10607
rect 0 10065 5573 10075
rect 0 9519 577836 10065
rect 0 9509 30045 9519
rect 0 8977 10265 8987
rect 0 8431 577836 8977
rect 0 8421 48353 8431
rect 0 7889 10081 7899
rect 0 7343 577836 7889
rect 0 7333 4561 7343
rect 0 6801 12473 6811
rect 0 6255 577836 6801
rect 0 6245 17349 6255
rect 0 5713 36853 5723
rect 0 5167 577836 5713
rect 0 5157 63993 5167
rect 0 4625 8793 4635
rect 0 4079 577836 4625
rect 0 4069 26641 4079
rect 0 3537 12749 3547
rect 0 2991 577836 3537
rect 0 2981 5941 2991
rect 0 2449 68777 2459
rect 0 2138 577836 2449
<< obsli1 >>
rect 38 765 577798 119731
<< obsm1 >>
rect 38 8 577798 120012
<< metal2 >>
rect 884 0 940 800
rect 4748 0 4804 800
rect 8704 0 8760 800
rect 12660 0 12716 800
rect 16616 0 16672 800
rect 20572 0 20628 800
rect 24528 0 24584 800
rect 28484 0 28540 800
rect 32440 0 32496 800
rect 36304 0 36360 800
rect 40260 0 40316 800
rect 44216 0 44272 800
rect 48172 0 48228 800
rect 52128 0 52184 800
rect 56084 0 56140 800
rect 60040 0 60096 800
rect 63996 0 64052 800
rect 67952 0 68008 800
rect 71816 0 71872 800
rect 75772 0 75828 800
rect 79728 0 79784 800
rect 83684 0 83740 800
rect 87640 0 87696 800
rect 91596 0 91652 800
rect 95552 0 95608 800
rect 99508 0 99564 800
rect 103372 0 103428 800
rect 107328 0 107384 800
rect 111284 0 111340 800
rect 115240 0 115296 800
rect 119196 0 119252 800
rect 123152 0 123208 800
rect 127108 0 127164 800
rect 131064 0 131120 800
rect 135020 0 135076 800
rect 138884 0 138940 800
rect 142840 0 142896 800
rect 146796 0 146852 800
rect 150752 0 150808 800
rect 154708 0 154764 800
rect 158664 0 158720 800
rect 162620 0 162676 800
rect 166576 0 166632 800
rect 170532 0 170588 800
rect 174396 0 174452 800
rect 178352 0 178408 800
rect 182308 0 182364 800
rect 186264 0 186320 800
rect 190220 0 190276 800
rect 194176 0 194232 800
rect 198132 0 198188 800
rect 202088 0 202144 800
rect 205952 0 206008 800
rect 209908 0 209964 800
rect 213864 0 213920 800
rect 217820 0 217876 800
rect 221776 0 221832 800
rect 225732 0 225788 800
rect 229688 0 229744 800
rect 233644 0 233700 800
rect 237600 0 237656 800
rect 241464 0 241520 800
rect 245420 0 245476 800
rect 249376 0 249432 800
rect 253332 0 253388 800
rect 257288 0 257344 800
rect 261244 0 261300 800
rect 265200 0 265256 800
rect 269156 0 269212 800
rect 273112 0 273168 800
rect 276976 0 277032 800
rect 280932 0 280988 800
rect 284888 0 284944 800
rect 288844 0 288900 800
rect 292800 0 292856 800
rect 296756 0 296812 800
rect 300712 0 300768 800
rect 304668 0 304724 800
rect 308532 0 308588 800
rect 312488 0 312544 800
rect 316444 0 316500 800
rect 320400 0 320456 800
rect 324356 0 324412 800
rect 328312 0 328368 800
rect 332268 0 332324 800
rect 336224 0 336280 800
rect 340180 0 340236 800
rect 344044 0 344100 800
rect 348000 0 348056 800
rect 351956 0 352012 800
rect 355912 0 355968 800
rect 359868 0 359924 800
rect 363824 0 363880 800
rect 367780 0 367836 800
rect 371736 0 371792 800
rect 375692 0 375748 800
rect 379556 0 379612 800
rect 383512 0 383568 800
rect 387468 0 387524 800
rect 391424 0 391480 800
rect 395380 0 395436 800
rect 399336 0 399392 800
rect 403292 0 403348 800
rect 407248 0 407304 800
rect 411112 0 411168 800
rect 415068 0 415124 800
rect 419024 0 419080 800
rect 422980 0 423036 800
rect 426936 0 426992 800
rect 430892 0 430948 800
rect 434848 0 434904 800
rect 438804 0 438860 800
rect 442760 0 442816 800
rect 446624 0 446680 800
rect 450580 0 450636 800
rect 454536 0 454592 800
rect 458492 0 458548 800
rect 462448 0 462504 800
rect 466404 0 466460 800
rect 470360 0 470416 800
rect 474316 0 474372 800
rect 478272 0 478328 800
rect 482136 0 482192 800
rect 486092 0 486148 800
rect 490048 0 490104 800
rect 494004 0 494060 800
rect 497960 0 498016 800
rect 501916 0 501972 800
rect 505872 0 505928 800
rect 509828 0 509884 800
rect 513692 0 513748 800
rect 517648 0 517704 800
rect 521604 0 521660 800
rect 525560 0 525616 800
rect 529516 0 529572 800
rect 533472 0 533528 800
rect 537428 0 537484 800
rect 541384 0 541440 800
rect 545340 0 545396 800
rect 549204 0 549260 800
rect 553160 0 553216 800
rect 557116 0 557172 800
rect 561072 0 561128 800
rect 565028 0 565084 800
rect 568984 0 569040 800
rect 572940 0 572996 800
rect 576896 0 576952 800
<< obsm2 >>
rect 426 856 577410 120018
rect 426 2 828 856
rect 996 2 4692 856
rect 4860 2 8648 856
rect 8816 2 12604 856
rect 12772 2 16560 856
rect 16728 2 20516 856
rect 20684 2 24472 856
rect 24640 2 28428 856
rect 28596 2 32384 856
rect 32552 2 36248 856
rect 36416 2 40204 856
rect 40372 2 44160 856
rect 44328 2 48116 856
rect 48284 2 52072 856
rect 52240 2 56028 856
rect 56196 2 59984 856
rect 60152 2 63940 856
rect 64108 2 67896 856
rect 68064 2 71760 856
rect 71928 2 75716 856
rect 75884 2 79672 856
rect 79840 2 83628 856
rect 83796 2 87584 856
rect 87752 2 91540 856
rect 91708 2 95496 856
rect 95664 2 99452 856
rect 99620 2 103316 856
rect 103484 2 107272 856
rect 107440 2 111228 856
rect 111396 2 115184 856
rect 115352 2 119140 856
rect 119308 2 123096 856
rect 123264 2 127052 856
rect 127220 2 131008 856
rect 131176 2 134964 856
rect 135132 2 138828 856
rect 138996 2 142784 856
rect 142952 2 146740 856
rect 146908 2 150696 856
rect 150864 2 154652 856
rect 154820 2 158608 856
rect 158776 2 162564 856
rect 162732 2 166520 856
rect 166688 2 170476 856
rect 170644 2 174340 856
rect 174508 2 178296 856
rect 178464 2 182252 856
rect 182420 2 186208 856
rect 186376 2 190164 856
rect 190332 2 194120 856
rect 194288 2 198076 856
rect 198244 2 202032 856
rect 202200 2 205896 856
rect 206064 2 209852 856
rect 210020 2 213808 856
rect 213976 2 217764 856
rect 217932 2 221720 856
rect 221888 2 225676 856
rect 225844 2 229632 856
rect 229800 2 233588 856
rect 233756 2 237544 856
rect 237712 2 241408 856
rect 241576 2 245364 856
rect 245532 2 249320 856
rect 249488 2 253276 856
rect 253444 2 257232 856
rect 257400 2 261188 856
rect 261356 2 265144 856
rect 265312 2 269100 856
rect 269268 2 273056 856
rect 273224 2 276920 856
rect 277088 2 280876 856
rect 281044 2 284832 856
rect 285000 2 288788 856
rect 288956 2 292744 856
rect 292912 2 296700 856
rect 296868 2 300656 856
rect 300824 2 304612 856
rect 304780 2 308476 856
rect 308644 2 312432 856
rect 312600 2 316388 856
rect 316556 2 320344 856
rect 320512 2 324300 856
rect 324468 2 328256 856
rect 328424 2 332212 856
rect 332380 2 336168 856
rect 336336 2 340124 856
rect 340292 2 343988 856
rect 344156 2 347944 856
rect 348112 2 351900 856
rect 352068 2 355856 856
rect 356024 2 359812 856
rect 359980 2 363768 856
rect 363936 2 367724 856
rect 367892 2 371680 856
rect 371848 2 375636 856
rect 375804 2 379500 856
rect 379668 2 383456 856
rect 383624 2 387412 856
rect 387580 2 391368 856
rect 391536 2 395324 856
rect 395492 2 399280 856
rect 399448 2 403236 856
rect 403404 2 407192 856
rect 407360 2 411056 856
rect 411224 2 415012 856
rect 415180 2 418968 856
rect 419136 2 422924 856
rect 423092 2 426880 856
rect 427048 2 430836 856
rect 431004 2 434792 856
rect 434960 2 438748 856
rect 438916 2 442704 856
rect 442872 2 446568 856
rect 446736 2 450524 856
rect 450692 2 454480 856
rect 454648 2 458436 856
rect 458604 2 462392 856
rect 462560 2 466348 856
rect 466516 2 470304 856
rect 470472 2 474260 856
rect 474428 2 478216 856
rect 478384 2 482080 856
rect 482248 2 486036 856
rect 486204 2 489992 856
rect 490160 2 493948 856
rect 494116 2 497904 856
rect 498072 2 501860 856
rect 502028 2 505816 856
rect 505984 2 509772 856
rect 509940 2 513636 856
rect 513804 2 517592 856
rect 517760 2 521548 856
rect 521716 2 525504 856
rect 525672 2 529460 856
rect 529628 2 533416 856
rect 533584 2 537372 856
rect 537540 2 541328 856
rect 541496 2 545284 856
rect 545452 2 549148 856
rect 549316 2 553104 856
rect 553272 2 557060 856
rect 557228 2 561016 856
rect 561184 2 564972 856
rect 565140 2 568928 856
rect 569096 2 572884 856
rect 573052 2 576840 856
rect 577008 2 577410 856
<< obsm3 >>
rect 511 35 577233 119917
<< metal4 >>
rect 3142 2128 3462 117552
rect 3802 2176 4122 117504
rect 4462 2176 4782 117504
rect 5122 2176 5442 117504
rect 18502 2128 18822 117552
rect 19162 2176 19482 117504
rect 19822 2176 20142 117504
rect 20482 2176 20802 117504
rect 33862 2128 34182 117552
rect 34522 2176 34842 117504
rect 35182 2176 35502 117504
rect 35842 2176 36162 117504
rect 49222 2128 49542 117552
rect 49882 2176 50202 117504
rect 50542 2176 50862 117504
rect 51202 2176 51522 117504
rect 64582 2128 64902 117552
rect 65242 2176 65562 117504
rect 65902 2176 66222 117504
rect 66562 2176 66882 117504
rect 79942 2128 80262 117552
rect 80602 2176 80922 117504
rect 81262 2176 81582 117504
rect 81922 2176 82242 117504
rect 95302 2128 95622 117552
rect 95962 2176 96282 117504
rect 96622 2176 96942 117504
rect 97282 2176 97602 117504
rect 110662 2128 110982 117552
rect 111322 2176 111642 117504
rect 111982 2176 112302 117504
rect 112642 2176 112962 117504
rect 126022 2128 126342 117552
rect 126682 2176 127002 117504
rect 127342 2176 127662 117504
rect 128002 2176 128322 117504
rect 141382 2128 141702 117552
rect 142042 2176 142362 117504
rect 142702 2176 143022 117504
rect 143362 2176 143682 117504
rect 156742 2128 157062 117552
rect 157402 2176 157722 117504
rect 158062 2176 158382 117504
rect 158722 2176 159042 117504
rect 172102 2128 172422 117552
rect 172762 2176 173082 117504
rect 173422 2176 173742 117504
rect 174082 2176 174402 117504
rect 187462 2128 187782 117552
rect 188122 2176 188442 117504
rect 188782 2176 189102 117504
rect 189442 2176 189762 117504
rect 202822 2128 203142 117552
rect 203482 2176 203802 117504
rect 204142 2176 204462 117504
rect 204802 2176 205122 117504
rect 218182 2128 218502 117552
rect 218842 2176 219162 117504
rect 219502 2176 219822 117504
rect 220162 2176 220482 117504
rect 233542 2128 233862 117552
rect 234202 2176 234522 117504
rect 234862 2176 235182 117504
rect 235522 2176 235842 117504
rect 248902 2128 249222 117552
rect 249562 2176 249882 117504
rect 250222 2176 250542 117504
rect 250882 2176 251202 117504
rect 264262 2128 264582 117552
rect 264922 2176 265242 117504
rect 265582 2176 265902 117504
rect 266242 2176 266562 117504
rect 279622 2128 279942 117552
rect 280282 2176 280602 117504
rect 280942 2176 281262 117504
rect 281602 2176 281922 117504
rect 294982 2128 295302 117552
rect 295642 2176 295962 117504
rect 296302 2176 296622 117504
rect 296962 2176 297282 117504
rect 310342 2128 310662 117552
rect 311002 2176 311322 117504
rect 311662 2176 311982 117504
rect 312322 2176 312642 117504
rect 325702 2128 326022 117552
rect 326362 2176 326682 117504
rect 327022 2176 327342 117504
rect 327682 2176 328002 117504
rect 341062 2128 341382 117552
rect 341722 2176 342042 117504
rect 342382 2176 342702 117504
rect 343042 2176 343362 117504
rect 356422 2128 356742 117552
rect 357082 2176 357402 117504
rect 357742 2176 358062 117504
rect 358402 2176 358722 117504
rect 371782 2128 372102 117552
rect 372442 2176 372762 117504
rect 373102 2176 373422 117504
rect 373762 2176 374082 117504
rect 387142 2128 387462 117552
rect 387802 2176 388122 117504
rect 388462 2176 388782 117504
rect 389122 2176 389442 117504
rect 402502 2128 402822 117552
rect 403162 2176 403482 117504
rect 403822 2176 404142 117504
rect 404482 2176 404802 117504
rect 417862 2128 418182 117552
rect 418522 2176 418842 117504
rect 419182 2176 419502 117504
rect 419842 2176 420162 117504
rect 433222 2128 433542 117552
rect 433882 2176 434202 117504
rect 434542 2176 434862 117504
rect 435202 2176 435522 117504
rect 448582 2128 448902 117552
rect 449242 2176 449562 117504
rect 449902 2176 450222 117504
rect 450562 2176 450882 117504
rect 463942 2128 464262 117552
rect 464602 2176 464922 117504
rect 465262 2176 465582 117504
rect 465922 2176 466242 117504
rect 479302 2128 479622 117552
rect 479962 2176 480282 117504
rect 480622 2176 480942 117504
rect 481282 2176 481602 117504
rect 494662 2128 494982 117552
rect 495322 2176 495642 117504
rect 495982 2176 496302 117504
rect 496642 2176 496962 117504
rect 510022 2128 510342 117552
rect 510682 2176 511002 117504
rect 511342 2176 511662 117504
rect 512002 2176 512322 117504
rect 525382 2128 525702 117552
rect 526042 2176 526362 117504
rect 526702 2176 527022 117504
rect 527362 2176 527682 117504
rect 540742 2128 541062 117552
rect 541402 2176 541722 117504
rect 542062 2176 542382 117504
rect 542722 2176 543042 117504
rect 556102 2128 556422 117552
rect 556762 2176 557082 117504
rect 557422 2176 557742 117504
rect 558082 2176 558402 117504
rect 571462 2128 571782 117552
rect 572122 2176 572442 117504
rect 572782 2176 573102 117504
rect 573442 2176 573762 117504
<< obsm4 >>
rect 18313 117632 559339 119917
rect 18313 2048 18422 117632
rect 18902 117584 33782 117632
rect 18902 2096 19082 117584
rect 19562 2096 19742 117584
rect 20222 2096 20402 117584
rect 20882 2096 33782 117584
rect 34262 117584 49142 117632
rect 18902 2048 33782 2096
rect 34262 2096 34442 117584
rect 34922 2096 35102 117584
rect 35582 2096 35762 117584
rect 36242 2096 49142 117584
rect 49622 117584 64502 117632
rect 34262 2048 49142 2096
rect 49622 2096 49802 117584
rect 50282 2096 50462 117584
rect 50942 2096 51122 117584
rect 51602 2096 64502 117584
rect 64982 117584 79862 117632
rect 49622 2048 64502 2096
rect 64982 2096 65162 117584
rect 65642 2096 65822 117584
rect 66302 2096 66482 117584
rect 66962 2096 79862 117584
rect 80342 117584 95222 117632
rect 64982 2048 79862 2096
rect 80342 2096 80522 117584
rect 81002 2096 81182 117584
rect 81662 2096 81842 117584
rect 82322 2096 95222 117584
rect 95702 117584 110582 117632
rect 80342 2048 95222 2096
rect 95702 2096 95882 117584
rect 96362 2096 96542 117584
rect 97022 2096 97202 117584
rect 97682 2096 110582 117584
rect 111062 117584 125942 117632
rect 95702 2048 110582 2096
rect 111062 2096 111242 117584
rect 111722 2096 111902 117584
rect 112382 2096 112562 117584
rect 113042 2096 125942 117584
rect 126422 117584 141302 117632
rect 111062 2048 125942 2096
rect 126422 2096 126602 117584
rect 127082 2096 127262 117584
rect 127742 2096 127922 117584
rect 128402 2096 141302 117584
rect 141782 117584 156662 117632
rect 126422 2048 141302 2096
rect 141782 2096 141962 117584
rect 142442 2096 142622 117584
rect 143102 2096 143282 117584
rect 143762 2096 156662 117584
rect 157142 117584 172022 117632
rect 141782 2048 156662 2096
rect 157142 2096 157322 117584
rect 157802 2096 157982 117584
rect 158462 2096 158642 117584
rect 159122 2096 172022 117584
rect 172502 117584 187382 117632
rect 157142 2048 172022 2096
rect 172502 2096 172682 117584
rect 173162 2096 173342 117584
rect 173822 2096 174002 117584
rect 174482 2096 187382 117584
rect 187862 117584 202742 117632
rect 172502 2048 187382 2096
rect 187862 2096 188042 117584
rect 188522 2096 188702 117584
rect 189182 2096 189362 117584
rect 189842 2096 202742 117584
rect 203222 117584 218102 117632
rect 187862 2048 202742 2096
rect 203222 2096 203402 117584
rect 203882 2096 204062 117584
rect 204542 2096 204722 117584
rect 205202 2096 218102 117584
rect 218582 117584 233462 117632
rect 203222 2048 218102 2096
rect 218582 2096 218762 117584
rect 219242 2096 219422 117584
rect 219902 2096 220082 117584
rect 220562 2096 233462 117584
rect 233942 117584 248822 117632
rect 218582 2048 233462 2096
rect 233942 2096 234122 117584
rect 234602 2096 234782 117584
rect 235262 2096 235442 117584
rect 235922 2096 248822 117584
rect 249302 117584 264182 117632
rect 233942 2048 248822 2096
rect 249302 2096 249482 117584
rect 249962 2096 250142 117584
rect 250622 2096 250802 117584
rect 251282 2096 264182 117584
rect 264662 117584 279542 117632
rect 249302 2048 264182 2096
rect 264662 2096 264842 117584
rect 265322 2096 265502 117584
rect 265982 2096 266162 117584
rect 266642 2096 279542 117584
rect 280022 117584 294902 117632
rect 264662 2048 279542 2096
rect 280022 2096 280202 117584
rect 280682 2096 280862 117584
rect 281342 2096 281522 117584
rect 282002 2096 294902 117584
rect 295382 117584 310262 117632
rect 280022 2048 294902 2096
rect 295382 2096 295562 117584
rect 296042 2096 296222 117584
rect 296702 2096 296882 117584
rect 297362 2096 310262 117584
rect 310742 117584 325622 117632
rect 295382 2048 310262 2096
rect 310742 2096 310922 117584
rect 311402 2096 311582 117584
rect 312062 2096 312242 117584
rect 312722 2096 325622 117584
rect 326102 117584 340982 117632
rect 310742 2048 325622 2096
rect 326102 2096 326282 117584
rect 326762 2096 326942 117584
rect 327422 2096 327602 117584
rect 328082 2096 340982 117584
rect 341462 117584 356342 117632
rect 326102 2048 340982 2096
rect 341462 2096 341642 117584
rect 342122 2096 342302 117584
rect 342782 2096 342962 117584
rect 343442 2096 356342 117584
rect 356822 117584 371702 117632
rect 341462 2048 356342 2096
rect 356822 2096 357002 117584
rect 357482 2096 357662 117584
rect 358142 2096 358322 117584
rect 358802 2096 371702 117584
rect 372182 117584 387062 117632
rect 356822 2048 371702 2096
rect 372182 2096 372362 117584
rect 372842 2096 373022 117584
rect 373502 2096 373682 117584
rect 374162 2096 387062 117584
rect 387542 117584 402422 117632
rect 372182 2048 387062 2096
rect 387542 2096 387722 117584
rect 388202 2096 388382 117584
rect 388862 2096 389042 117584
rect 389522 2096 402422 117584
rect 402902 117584 417782 117632
rect 387542 2048 402422 2096
rect 402902 2096 403082 117584
rect 403562 2096 403742 117584
rect 404222 2096 404402 117584
rect 404882 2096 417782 117584
rect 418262 117584 433142 117632
rect 402902 2048 417782 2096
rect 418262 2096 418442 117584
rect 418922 2096 419102 117584
rect 419582 2096 419762 117584
rect 420242 2096 433142 117584
rect 433622 117584 448502 117632
rect 418262 2048 433142 2096
rect 433622 2096 433802 117584
rect 434282 2096 434462 117584
rect 434942 2096 435122 117584
rect 435602 2096 448502 117584
rect 448982 117584 463862 117632
rect 433622 2048 448502 2096
rect 448982 2096 449162 117584
rect 449642 2096 449822 117584
rect 450302 2096 450482 117584
rect 450962 2096 463862 117584
rect 464342 117584 479222 117632
rect 448982 2048 463862 2096
rect 464342 2096 464522 117584
rect 465002 2096 465182 117584
rect 465662 2096 465842 117584
rect 466322 2096 479222 117584
rect 479702 117584 494582 117632
rect 464342 2048 479222 2096
rect 479702 2096 479882 117584
rect 480362 2096 480542 117584
rect 481022 2096 481202 117584
rect 481682 2096 494582 117584
rect 495062 117584 509942 117632
rect 479702 2048 494582 2096
rect 495062 2096 495242 117584
rect 495722 2096 495902 117584
rect 496382 2096 496562 117584
rect 497042 2096 509942 117584
rect 510422 117584 525302 117632
rect 495062 2048 509942 2096
rect 510422 2096 510602 117584
rect 511082 2096 511262 117584
rect 511742 2096 511922 117584
rect 512402 2096 525302 117584
rect 525782 117584 540662 117632
rect 510422 2048 525302 2096
rect 525782 2096 525962 117584
rect 526442 2096 526622 117584
rect 527102 2096 527282 117584
rect 527762 2096 540662 117584
rect 541142 117584 556022 117632
rect 525782 2048 540662 2096
rect 541142 2096 541322 117584
rect 541802 2096 541982 117584
rect 542462 2096 542642 117584
rect 543122 2096 556022 117584
rect 556502 117584 559339 117632
rect 541142 2048 556022 2096
rect 556502 2096 556682 117584
rect 557162 2096 557342 117584
rect 557822 2096 558002 117584
rect 558482 2096 559339 117584
rect 556502 2048 559339 2096
rect 18313 35 559339 2048
<< labels >>
rlabel metal2 s 505872 0 505928 800 6 A[0]
port 1 nsew signal input
rlabel metal2 s 509828 0 509884 800 6 A[1]
port 2 nsew signal input
rlabel metal2 s 513692 0 513748 800 6 A[2]
port 3 nsew signal input
rlabel metal2 s 517648 0 517704 800 6 A[3]
port 4 nsew signal input
rlabel metal2 s 521604 0 521660 800 6 A[4]
port 5 nsew signal input
rlabel metal2 s 525560 0 525616 800 6 A[5]
port 6 nsew signal input
rlabel metal2 s 529516 0 529572 800 6 A[6]
port 7 nsew signal input
rlabel metal2 s 533472 0 533528 800 6 A[7]
port 8 nsew signal input
rlabel metal2 s 537428 0 537484 800 6 A[8]
port 9 nsew signal input
rlabel metal2 s 541384 0 541440 800 6 CLK
port 10 nsew signal input
rlabel metal2 s 253332 0 253388 800 6 Di[0]
port 11 nsew signal input
rlabel metal2 s 292800 0 292856 800 6 Di[10]
port 12 nsew signal input
rlabel metal2 s 296756 0 296812 800 6 Di[11]
port 13 nsew signal input
rlabel metal2 s 300712 0 300768 800 6 Di[12]
port 14 nsew signal input
rlabel metal2 s 304668 0 304724 800 6 Di[13]
port 15 nsew signal input
rlabel metal2 s 308532 0 308588 800 6 Di[14]
port 16 nsew signal input
rlabel metal2 s 312488 0 312544 800 6 Di[15]
port 17 nsew signal input
rlabel metal2 s 316444 0 316500 800 6 Di[16]
port 18 nsew signal input
rlabel metal2 s 320400 0 320456 800 6 Di[17]
port 19 nsew signal input
rlabel metal2 s 324356 0 324412 800 6 Di[18]
port 20 nsew signal input
rlabel metal2 s 328312 0 328368 800 6 Di[19]
port 21 nsew signal input
rlabel metal2 s 257288 0 257344 800 6 Di[1]
port 22 nsew signal input
rlabel metal2 s 332268 0 332324 800 6 Di[20]
port 23 nsew signal input
rlabel metal2 s 336224 0 336280 800 6 Di[21]
port 24 nsew signal input
rlabel metal2 s 340180 0 340236 800 6 Di[22]
port 25 nsew signal input
rlabel metal2 s 344044 0 344100 800 6 Di[23]
port 26 nsew signal input
rlabel metal2 s 348000 0 348056 800 6 Di[24]
port 27 nsew signal input
rlabel metal2 s 351956 0 352012 800 6 Di[25]
port 28 nsew signal input
rlabel metal2 s 355912 0 355968 800 6 Di[26]
port 29 nsew signal input
rlabel metal2 s 359868 0 359924 800 6 Di[27]
port 30 nsew signal input
rlabel metal2 s 363824 0 363880 800 6 Di[28]
port 31 nsew signal input
rlabel metal2 s 367780 0 367836 800 6 Di[29]
port 32 nsew signal input
rlabel metal2 s 261244 0 261300 800 6 Di[2]
port 33 nsew signal input
rlabel metal2 s 371736 0 371792 800 6 Di[30]
port 34 nsew signal input
rlabel metal2 s 375692 0 375748 800 6 Di[31]
port 35 nsew signal input
rlabel metal2 s 379556 0 379612 800 6 Di[32]
port 36 nsew signal input
rlabel metal2 s 383512 0 383568 800 6 Di[33]
port 37 nsew signal input
rlabel metal2 s 387468 0 387524 800 6 Di[34]
port 38 nsew signal input
rlabel metal2 s 391424 0 391480 800 6 Di[35]
port 39 nsew signal input
rlabel metal2 s 395380 0 395436 800 6 Di[36]
port 40 nsew signal input
rlabel metal2 s 399336 0 399392 800 6 Di[37]
port 41 nsew signal input
rlabel metal2 s 403292 0 403348 800 6 Di[38]
port 42 nsew signal input
rlabel metal2 s 407248 0 407304 800 6 Di[39]
port 43 nsew signal input
rlabel metal2 s 265200 0 265256 800 6 Di[3]
port 44 nsew signal input
rlabel metal2 s 411112 0 411168 800 6 Di[40]
port 45 nsew signal input
rlabel metal2 s 415068 0 415124 800 6 Di[41]
port 46 nsew signal input
rlabel metal2 s 419024 0 419080 800 6 Di[42]
port 47 nsew signal input
rlabel metal2 s 422980 0 423036 800 6 Di[43]
port 48 nsew signal input
rlabel metal2 s 426936 0 426992 800 6 Di[44]
port 49 nsew signal input
rlabel metal2 s 430892 0 430948 800 6 Di[45]
port 50 nsew signal input
rlabel metal2 s 434848 0 434904 800 6 Di[46]
port 51 nsew signal input
rlabel metal2 s 438804 0 438860 800 6 Di[47]
port 52 nsew signal input
rlabel metal2 s 442760 0 442816 800 6 Di[48]
port 53 nsew signal input
rlabel metal2 s 446624 0 446680 800 6 Di[49]
port 54 nsew signal input
rlabel metal2 s 269156 0 269212 800 6 Di[4]
port 55 nsew signal input
rlabel metal2 s 450580 0 450636 800 6 Di[50]
port 56 nsew signal input
rlabel metal2 s 454536 0 454592 800 6 Di[51]
port 57 nsew signal input
rlabel metal2 s 458492 0 458548 800 6 Di[52]
port 58 nsew signal input
rlabel metal2 s 462448 0 462504 800 6 Di[53]
port 59 nsew signal input
rlabel metal2 s 466404 0 466460 800 6 Di[54]
port 60 nsew signal input
rlabel metal2 s 470360 0 470416 800 6 Di[55]
port 61 nsew signal input
rlabel metal2 s 474316 0 474372 800 6 Di[56]
port 62 nsew signal input
rlabel metal2 s 478272 0 478328 800 6 Di[57]
port 63 nsew signal input
rlabel metal2 s 482136 0 482192 800 6 Di[58]
port 64 nsew signal input
rlabel metal2 s 486092 0 486148 800 6 Di[59]
port 65 nsew signal input
rlabel metal2 s 273112 0 273168 800 6 Di[5]
port 66 nsew signal input
rlabel metal2 s 490048 0 490104 800 6 Di[60]
port 67 nsew signal input
rlabel metal2 s 494004 0 494060 800 6 Di[61]
port 68 nsew signal input
rlabel metal2 s 497960 0 498016 800 6 Di[62]
port 69 nsew signal input
rlabel metal2 s 501916 0 501972 800 6 Di[63]
port 70 nsew signal input
rlabel metal2 s 276976 0 277032 800 6 Di[6]
port 71 nsew signal input
rlabel metal2 s 280932 0 280988 800 6 Di[7]
port 72 nsew signal input
rlabel metal2 s 284888 0 284944 800 6 Di[8]
port 73 nsew signal input
rlabel metal2 s 288844 0 288900 800 6 Di[9]
port 74 nsew signal input
rlabel metal2 s 884 0 940 800 6 Do[0]
port 75 nsew signal output
rlabel metal2 s 40260 0 40316 800 6 Do[10]
port 76 nsew signal output
rlabel metal2 s 44216 0 44272 800 6 Do[11]
port 77 nsew signal output
rlabel metal2 s 48172 0 48228 800 6 Do[12]
port 78 nsew signal output
rlabel metal2 s 52128 0 52184 800 6 Do[13]
port 79 nsew signal output
rlabel metal2 s 56084 0 56140 800 6 Do[14]
port 80 nsew signal output
rlabel metal2 s 60040 0 60096 800 6 Do[15]
port 81 nsew signal output
rlabel metal2 s 63996 0 64052 800 6 Do[16]
port 82 nsew signal output
rlabel metal2 s 67952 0 68008 800 6 Do[17]
port 83 nsew signal output
rlabel metal2 s 71816 0 71872 800 6 Do[18]
port 84 nsew signal output
rlabel metal2 s 75772 0 75828 800 6 Do[19]
port 85 nsew signal output
rlabel metal2 s 4748 0 4804 800 6 Do[1]
port 86 nsew signal output
rlabel metal2 s 79728 0 79784 800 6 Do[20]
port 87 nsew signal output
rlabel metal2 s 83684 0 83740 800 6 Do[21]
port 88 nsew signal output
rlabel metal2 s 87640 0 87696 800 6 Do[22]
port 89 nsew signal output
rlabel metal2 s 91596 0 91652 800 6 Do[23]
port 90 nsew signal output
rlabel metal2 s 95552 0 95608 800 6 Do[24]
port 91 nsew signal output
rlabel metal2 s 99508 0 99564 800 6 Do[25]
port 92 nsew signal output
rlabel metal2 s 103372 0 103428 800 6 Do[26]
port 93 nsew signal output
rlabel metal2 s 107328 0 107384 800 6 Do[27]
port 94 nsew signal output
rlabel metal2 s 111284 0 111340 800 6 Do[28]
port 95 nsew signal output
rlabel metal2 s 115240 0 115296 800 6 Do[29]
port 96 nsew signal output
rlabel metal2 s 8704 0 8760 800 6 Do[2]
port 97 nsew signal output
rlabel metal2 s 119196 0 119252 800 6 Do[30]
port 98 nsew signal output
rlabel metal2 s 123152 0 123208 800 6 Do[31]
port 99 nsew signal output
rlabel metal2 s 127108 0 127164 800 6 Do[32]
port 100 nsew signal output
rlabel metal2 s 131064 0 131120 800 6 Do[33]
port 101 nsew signal output
rlabel metal2 s 135020 0 135076 800 6 Do[34]
port 102 nsew signal output
rlabel metal2 s 138884 0 138940 800 6 Do[35]
port 103 nsew signal output
rlabel metal2 s 142840 0 142896 800 6 Do[36]
port 104 nsew signal output
rlabel metal2 s 146796 0 146852 800 6 Do[37]
port 105 nsew signal output
rlabel metal2 s 150752 0 150808 800 6 Do[38]
port 106 nsew signal output
rlabel metal2 s 154708 0 154764 800 6 Do[39]
port 107 nsew signal output
rlabel metal2 s 12660 0 12716 800 6 Do[3]
port 108 nsew signal output
rlabel metal2 s 158664 0 158720 800 6 Do[40]
port 109 nsew signal output
rlabel metal2 s 162620 0 162676 800 6 Do[41]
port 110 nsew signal output
rlabel metal2 s 166576 0 166632 800 6 Do[42]
port 111 nsew signal output
rlabel metal2 s 170532 0 170588 800 6 Do[43]
port 112 nsew signal output
rlabel metal2 s 174396 0 174452 800 6 Do[44]
port 113 nsew signal output
rlabel metal2 s 178352 0 178408 800 6 Do[45]
port 114 nsew signal output
rlabel metal2 s 182308 0 182364 800 6 Do[46]
port 115 nsew signal output
rlabel metal2 s 186264 0 186320 800 6 Do[47]
port 116 nsew signal output
rlabel metal2 s 190220 0 190276 800 6 Do[48]
port 117 nsew signal output
rlabel metal2 s 194176 0 194232 800 6 Do[49]
port 118 nsew signal output
rlabel metal2 s 16616 0 16672 800 6 Do[4]
port 119 nsew signal output
rlabel metal2 s 198132 0 198188 800 6 Do[50]
port 120 nsew signal output
rlabel metal2 s 202088 0 202144 800 6 Do[51]
port 121 nsew signal output
rlabel metal2 s 205952 0 206008 800 6 Do[52]
port 122 nsew signal output
rlabel metal2 s 209908 0 209964 800 6 Do[53]
port 123 nsew signal output
rlabel metal2 s 213864 0 213920 800 6 Do[54]
port 124 nsew signal output
rlabel metal2 s 217820 0 217876 800 6 Do[55]
port 125 nsew signal output
rlabel metal2 s 221776 0 221832 800 6 Do[56]
port 126 nsew signal output
rlabel metal2 s 225732 0 225788 800 6 Do[57]
port 127 nsew signal output
rlabel metal2 s 229688 0 229744 800 6 Do[58]
port 128 nsew signal output
rlabel metal2 s 233644 0 233700 800 6 Do[59]
port 129 nsew signal output
rlabel metal2 s 20572 0 20628 800 6 Do[5]
port 130 nsew signal output
rlabel metal2 s 237600 0 237656 800 6 Do[60]
port 131 nsew signal output
rlabel metal2 s 241464 0 241520 800 6 Do[61]
port 132 nsew signal output
rlabel metal2 s 245420 0 245476 800 6 Do[62]
port 133 nsew signal output
rlabel metal2 s 249376 0 249432 800 6 Do[63]
port 134 nsew signal output
rlabel metal2 s 24528 0 24584 800 6 Do[6]
port 135 nsew signal output
rlabel metal2 s 28484 0 28540 800 6 Do[7]
port 136 nsew signal output
rlabel metal2 s 32440 0 32496 800 6 Do[8]
port 137 nsew signal output
rlabel metal2 s 36304 0 36360 800 6 Do[9]
port 138 nsew signal output
rlabel metal2 s 576896 0 576952 800 6 EN
port 139 nsew signal input
rlabel metal2 s 545340 0 545396 800 6 WE[0]
port 140 nsew signal input
rlabel metal2 s 549204 0 549260 800 6 WE[1]
port 141 nsew signal input
rlabel metal2 s 553160 0 553216 800 6 WE[2]
port 142 nsew signal input
rlabel metal2 s 557116 0 557172 800 6 WE[3]
port 143 nsew signal input
rlabel metal2 s 561072 0 561128 800 6 WE[4]
port 144 nsew signal input
rlabel metal2 s 565028 0 565084 800 6 WE[5]
port 145 nsew signal input
rlabel metal2 s 568984 0 569040 800 6 WE[6]
port 146 nsew signal input
rlabel metal2 s 572940 0 572996 800 6 WE[7]
port 147 nsew signal input
rlabel metal4 s 556102 2128 556422 117552 6 vccd1
port 148 nsew power bidirectional
rlabel metal4 s 525382 2128 525702 117552 6 vccd1
port 149 nsew power bidirectional
rlabel metal4 s 494662 2128 494982 117552 6 vccd1
port 150 nsew power bidirectional
rlabel metal4 s 463942 2128 464262 117552 6 vccd1
port 151 nsew power bidirectional
rlabel metal4 s 433222 2128 433542 117552 6 vccd1
port 152 nsew power bidirectional
rlabel metal4 s 402502 2128 402822 117552 6 vccd1
port 153 nsew power bidirectional
rlabel metal4 s 371782 2128 372102 117552 6 vccd1
port 154 nsew power bidirectional
rlabel metal4 s 341062 2128 341382 117552 6 vccd1
port 155 nsew power bidirectional
rlabel metal4 s 310342 2128 310662 117552 6 vccd1
port 156 nsew power bidirectional
rlabel metal4 s 279622 2128 279942 117552 6 vccd1
port 157 nsew power bidirectional
rlabel metal4 s 248902 2128 249222 117552 6 vccd1
port 158 nsew power bidirectional
rlabel metal4 s 218182 2128 218502 117552 6 vccd1
port 159 nsew power bidirectional
rlabel metal4 s 187462 2128 187782 117552 6 vccd1
port 160 nsew power bidirectional
rlabel metal4 s 156742 2128 157062 117552 6 vccd1
port 161 nsew power bidirectional
rlabel metal4 s 126022 2128 126342 117552 6 vccd1
port 162 nsew power bidirectional
rlabel metal4 s 95302 2128 95622 117552 6 vccd1
port 163 nsew power bidirectional
rlabel metal4 s 64582 2128 64902 117552 6 vccd1
port 164 nsew power bidirectional
rlabel metal4 s 33862 2128 34182 117552 6 vccd1
port 165 nsew power bidirectional
rlabel metal4 s 3142 2128 3462 117552 6 vccd1
port 166 nsew power bidirectional
rlabel metal4 s 571462 2128 571782 117552 6 vssd1
port 167 nsew ground bidirectional
rlabel metal4 s 540742 2128 541062 117552 6 vssd1
port 168 nsew ground bidirectional
rlabel metal4 s 510022 2128 510342 117552 6 vssd1
port 169 nsew ground bidirectional
rlabel metal4 s 479302 2128 479622 117552 6 vssd1
port 170 nsew ground bidirectional
rlabel metal4 s 448582 2128 448902 117552 6 vssd1
port 171 nsew ground bidirectional
rlabel metal4 s 417862 2128 418182 117552 6 vssd1
port 172 nsew ground bidirectional
rlabel metal4 s 387142 2128 387462 117552 6 vssd1
port 173 nsew ground bidirectional
rlabel metal4 s 356422 2128 356742 117552 6 vssd1
port 174 nsew ground bidirectional
rlabel metal4 s 325702 2128 326022 117552 6 vssd1
port 175 nsew ground bidirectional
rlabel metal4 s 294982 2128 295302 117552 6 vssd1
port 176 nsew ground bidirectional
rlabel metal4 s 264262 2128 264582 117552 6 vssd1
port 177 nsew ground bidirectional
rlabel metal4 s 233542 2128 233862 117552 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 202822 2128 203142 117552 6 vssd1
port 179 nsew ground bidirectional
rlabel metal4 s 172102 2128 172422 117552 6 vssd1
port 180 nsew ground bidirectional
rlabel metal4 s 141382 2128 141702 117552 6 vssd1
port 181 nsew ground bidirectional
rlabel metal4 s 110662 2128 110982 117552 6 vssd1
port 182 nsew ground bidirectional
rlabel metal4 s 79942 2128 80262 117552 6 vssd1
port 183 nsew ground bidirectional
rlabel metal4 s 49222 2128 49542 117552 6 vssd1
port 184 nsew ground bidirectional
rlabel metal4 s 18502 2128 18822 117552 6 vssd1
port 185 nsew ground bidirectional
rlabel metal4 s 556762 2176 557082 117504 6 vccd2
port 186 nsew power bidirectional
rlabel metal4 s 526042 2176 526362 117504 6 vccd2
port 187 nsew power bidirectional
rlabel metal4 s 495322 2176 495642 117504 6 vccd2
port 188 nsew power bidirectional
rlabel metal4 s 464602 2176 464922 117504 6 vccd2
port 189 nsew power bidirectional
rlabel metal4 s 433882 2176 434202 117504 6 vccd2
port 190 nsew power bidirectional
rlabel metal4 s 403162 2176 403482 117504 6 vccd2
port 191 nsew power bidirectional
rlabel metal4 s 372442 2176 372762 117504 6 vccd2
port 192 nsew power bidirectional
rlabel metal4 s 341722 2176 342042 117504 6 vccd2
port 193 nsew power bidirectional
rlabel metal4 s 311002 2176 311322 117504 6 vccd2
port 194 nsew power bidirectional
rlabel metal4 s 280282 2176 280602 117504 6 vccd2
port 195 nsew power bidirectional
rlabel metal4 s 249562 2176 249882 117504 6 vccd2
port 196 nsew power bidirectional
rlabel metal4 s 218842 2176 219162 117504 6 vccd2
port 197 nsew power bidirectional
rlabel metal4 s 188122 2176 188442 117504 6 vccd2
port 198 nsew power bidirectional
rlabel metal4 s 157402 2176 157722 117504 6 vccd2
port 199 nsew power bidirectional
rlabel metal4 s 126682 2176 127002 117504 6 vccd2
port 200 nsew power bidirectional
rlabel metal4 s 95962 2176 96282 117504 6 vccd2
port 201 nsew power bidirectional
rlabel metal4 s 65242 2176 65562 117504 6 vccd2
port 202 nsew power bidirectional
rlabel metal4 s 34522 2176 34842 117504 6 vccd2
port 203 nsew power bidirectional
rlabel metal4 s 3802 2176 4122 117504 6 vccd2
port 204 nsew power bidirectional
rlabel metal4 s 572122 2176 572442 117504 6 vssd2
port 205 nsew ground bidirectional
rlabel metal4 s 541402 2176 541722 117504 6 vssd2
port 206 nsew ground bidirectional
rlabel metal4 s 510682 2176 511002 117504 6 vssd2
port 207 nsew ground bidirectional
rlabel metal4 s 479962 2176 480282 117504 6 vssd2
port 208 nsew ground bidirectional
rlabel metal4 s 449242 2176 449562 117504 6 vssd2
port 209 nsew ground bidirectional
rlabel metal4 s 418522 2176 418842 117504 6 vssd2
port 210 nsew ground bidirectional
rlabel metal4 s 387802 2176 388122 117504 6 vssd2
port 211 nsew ground bidirectional
rlabel metal4 s 357082 2176 357402 117504 6 vssd2
port 212 nsew ground bidirectional
rlabel metal4 s 326362 2176 326682 117504 6 vssd2
port 213 nsew ground bidirectional
rlabel metal4 s 295642 2176 295962 117504 6 vssd2
port 214 nsew ground bidirectional
rlabel metal4 s 264922 2176 265242 117504 6 vssd2
port 215 nsew ground bidirectional
rlabel metal4 s 234202 2176 234522 117504 6 vssd2
port 216 nsew ground bidirectional
rlabel metal4 s 203482 2176 203802 117504 6 vssd2
port 217 nsew ground bidirectional
rlabel metal4 s 172762 2176 173082 117504 6 vssd2
port 218 nsew ground bidirectional
rlabel metal4 s 142042 2176 142362 117504 6 vssd2
port 219 nsew ground bidirectional
rlabel metal4 s 111322 2176 111642 117504 6 vssd2
port 220 nsew ground bidirectional
rlabel metal4 s 80602 2176 80922 117504 6 vssd2
port 221 nsew ground bidirectional
rlabel metal4 s 49882 2176 50202 117504 6 vssd2
port 222 nsew ground bidirectional
rlabel metal4 s 19162 2176 19482 117504 6 vssd2
port 223 nsew ground bidirectional
rlabel metal4 s 557422 2176 557742 117504 6 vdda1
port 224 nsew power bidirectional
rlabel metal4 s 526702 2176 527022 117504 6 vdda1
port 225 nsew power bidirectional
rlabel metal4 s 495982 2176 496302 117504 6 vdda1
port 226 nsew power bidirectional
rlabel metal4 s 465262 2176 465582 117504 6 vdda1
port 227 nsew power bidirectional
rlabel metal4 s 434542 2176 434862 117504 6 vdda1
port 228 nsew power bidirectional
rlabel metal4 s 403822 2176 404142 117504 6 vdda1
port 229 nsew power bidirectional
rlabel metal4 s 373102 2176 373422 117504 6 vdda1
port 230 nsew power bidirectional
rlabel metal4 s 342382 2176 342702 117504 6 vdda1
port 231 nsew power bidirectional
rlabel metal4 s 311662 2176 311982 117504 6 vdda1
port 232 nsew power bidirectional
rlabel metal4 s 280942 2176 281262 117504 6 vdda1
port 233 nsew power bidirectional
rlabel metal4 s 250222 2176 250542 117504 6 vdda1
port 234 nsew power bidirectional
rlabel metal4 s 219502 2176 219822 117504 6 vdda1
port 235 nsew power bidirectional
rlabel metal4 s 188782 2176 189102 117504 6 vdda1
port 236 nsew power bidirectional
rlabel metal4 s 158062 2176 158382 117504 6 vdda1
port 237 nsew power bidirectional
rlabel metal4 s 127342 2176 127662 117504 6 vdda1
port 238 nsew power bidirectional
rlabel metal4 s 96622 2176 96942 117504 6 vdda1
port 239 nsew power bidirectional
rlabel metal4 s 65902 2176 66222 117504 6 vdda1
port 240 nsew power bidirectional
rlabel metal4 s 35182 2176 35502 117504 6 vdda1
port 241 nsew power bidirectional
rlabel metal4 s 4462 2176 4782 117504 6 vdda1
port 242 nsew power bidirectional
rlabel metal4 s 572782 2176 573102 117504 6 vssa1
port 243 nsew ground bidirectional
rlabel metal4 s 542062 2176 542382 117504 6 vssa1
port 244 nsew ground bidirectional
rlabel metal4 s 511342 2176 511662 117504 6 vssa1
port 245 nsew ground bidirectional
rlabel metal4 s 480622 2176 480942 117504 6 vssa1
port 246 nsew ground bidirectional
rlabel metal4 s 449902 2176 450222 117504 6 vssa1
port 247 nsew ground bidirectional
rlabel metal4 s 419182 2176 419502 117504 6 vssa1
port 248 nsew ground bidirectional
rlabel metal4 s 388462 2176 388782 117504 6 vssa1
port 249 nsew ground bidirectional
rlabel metal4 s 357742 2176 358062 117504 6 vssa1
port 250 nsew ground bidirectional
rlabel metal4 s 327022 2176 327342 117504 6 vssa1
port 251 nsew ground bidirectional
rlabel metal4 s 296302 2176 296622 117504 6 vssa1
port 252 nsew ground bidirectional
rlabel metal4 s 265582 2176 265902 117504 6 vssa1
port 253 nsew ground bidirectional
rlabel metal4 s 234862 2176 235182 117504 6 vssa1
port 254 nsew ground bidirectional
rlabel metal4 s 204142 2176 204462 117504 6 vssa1
port 255 nsew ground bidirectional
rlabel metal4 s 173422 2176 173742 117504 6 vssa1
port 256 nsew ground bidirectional
rlabel metal4 s 142702 2176 143022 117504 6 vssa1
port 257 nsew ground bidirectional
rlabel metal4 s 111982 2176 112302 117504 6 vssa1
port 258 nsew ground bidirectional
rlabel metal4 s 81262 2176 81582 117504 6 vssa1
port 259 nsew ground bidirectional
rlabel metal4 s 50542 2176 50862 117504 6 vssa1
port 260 nsew ground bidirectional
rlabel metal4 s 19822 2176 20142 117504 6 vssa1
port 261 nsew ground bidirectional
rlabel metal4 s 558082 2176 558402 117504 6 vdda2
port 262 nsew power bidirectional
rlabel metal4 s 527362 2176 527682 117504 6 vdda2
port 263 nsew power bidirectional
rlabel metal4 s 496642 2176 496962 117504 6 vdda2
port 264 nsew power bidirectional
rlabel metal4 s 465922 2176 466242 117504 6 vdda2
port 265 nsew power bidirectional
rlabel metal4 s 435202 2176 435522 117504 6 vdda2
port 266 nsew power bidirectional
rlabel metal4 s 404482 2176 404802 117504 6 vdda2
port 267 nsew power bidirectional
rlabel metal4 s 373762 2176 374082 117504 6 vdda2
port 268 nsew power bidirectional
rlabel metal4 s 343042 2176 343362 117504 6 vdda2
port 269 nsew power bidirectional
rlabel metal4 s 312322 2176 312642 117504 6 vdda2
port 270 nsew power bidirectional
rlabel metal4 s 281602 2176 281922 117504 6 vdda2
port 271 nsew power bidirectional
rlabel metal4 s 250882 2176 251202 117504 6 vdda2
port 272 nsew power bidirectional
rlabel metal4 s 220162 2176 220482 117504 6 vdda2
port 273 nsew power bidirectional
rlabel metal4 s 189442 2176 189762 117504 6 vdda2
port 274 nsew power bidirectional
rlabel metal4 s 158722 2176 159042 117504 6 vdda2
port 275 nsew power bidirectional
rlabel metal4 s 128002 2176 128322 117504 6 vdda2
port 276 nsew power bidirectional
rlabel metal4 s 97282 2176 97602 117504 6 vdda2
port 277 nsew power bidirectional
rlabel metal4 s 66562 2176 66882 117504 6 vdda2
port 278 nsew power bidirectional
rlabel metal4 s 35842 2176 36162 117504 6 vdda2
port 279 nsew power bidirectional
rlabel metal4 s 5122 2176 5442 117504 6 vdda2
port 280 nsew power bidirectional
rlabel metal4 s 573442 2176 573762 117504 6 vssa2
port 281 nsew ground bidirectional
rlabel metal4 s 542722 2176 543042 117504 6 vssa2
port 282 nsew ground bidirectional
rlabel metal4 s 512002 2176 512322 117504 6 vssa2
port 283 nsew ground bidirectional
rlabel metal4 s 481282 2176 481602 117504 6 vssa2
port 284 nsew ground bidirectional
rlabel metal4 s 450562 2176 450882 117504 6 vssa2
port 285 nsew ground bidirectional
rlabel metal4 s 419842 2176 420162 117504 6 vssa2
port 286 nsew ground bidirectional
rlabel metal4 s 389122 2176 389442 117504 6 vssa2
port 287 nsew ground bidirectional
rlabel metal4 s 358402 2176 358722 117504 6 vssa2
port 288 nsew ground bidirectional
rlabel metal4 s 327682 2176 328002 117504 6 vssa2
port 289 nsew ground bidirectional
rlabel metal4 s 296962 2176 297282 117504 6 vssa2
port 290 nsew ground bidirectional
rlabel metal4 s 266242 2176 266562 117504 6 vssa2
port 291 nsew ground bidirectional
rlabel metal4 s 235522 2176 235842 117504 6 vssa2
port 292 nsew ground bidirectional
rlabel metal4 s 204802 2176 205122 117504 6 vssa2
port 293 nsew ground bidirectional
rlabel metal4 s 174082 2176 174402 117504 6 vssa2
port 294 nsew ground bidirectional
rlabel metal4 s 143362 2176 143682 117504 6 vssa2
port 295 nsew ground bidirectional
rlabel metal4 s 112642 2176 112962 117504 6 vssa2
port 296 nsew ground bidirectional
rlabel metal4 s 81922 2176 82242 117504 6 vssa2
port 297 nsew ground bidirectional
rlabel metal4 s 51202 2176 51522 117504 6 vssa2
port 298 nsew ground bidirectional
rlabel metal4 s 20482 2176 20802 117504 6 vssa2
port 299 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 577836 120018
string LEFview TRUE
string GDS_FILE /project/openlane/RAM_512x64/runs/RAM_512x64/results/magic/RAM_512x64.gds
string GDS_END 236567988
string GDS_START 190756
<< end >>

