magic
tech sky130A
magscale 1 2
timestamp 1608847369
<< obsli1 >>
rect 38 1309 557742 157777
<< obsm1 >>
rect 38 1300 557742 157808
<< metal2 >>
rect 792 0 848 800
rect 4564 0 4620 800
rect 8336 0 8392 800
rect 12200 0 12256 800
rect 15972 0 16028 800
rect 19836 0 19892 800
rect 23608 0 23664 800
rect 27380 0 27436 800
rect 31244 0 31300 800
rect 35016 0 35072 800
rect 38880 0 38936 800
rect 42652 0 42708 800
rect 46424 0 46480 800
rect 50288 0 50344 800
rect 54060 0 54116 800
rect 57924 0 57980 800
rect 61696 0 61752 800
rect 65468 0 65524 800
rect 69332 0 69388 800
rect 73104 0 73160 800
rect 76968 0 77024 800
rect 80740 0 80796 800
rect 84512 0 84568 800
rect 88376 0 88432 800
rect 92148 0 92204 800
rect 96012 0 96068 800
rect 99784 0 99840 800
rect 103648 0 103704 800
rect 107420 0 107476 800
rect 111192 0 111248 800
rect 115056 0 115112 800
rect 118828 0 118884 800
rect 122692 0 122748 800
rect 126464 0 126520 800
rect 130236 0 130292 800
rect 134100 0 134156 800
rect 137872 0 137928 800
rect 141736 0 141792 800
rect 145508 0 145564 800
rect 149280 0 149336 800
rect 153144 0 153200 800
rect 156916 0 156972 800
rect 160780 0 160836 800
rect 164552 0 164608 800
rect 168324 0 168380 800
rect 172188 0 172244 800
rect 175960 0 176016 800
rect 179824 0 179880 800
rect 183596 0 183652 800
rect 187460 0 187516 800
rect 191232 0 191288 800
rect 195004 0 195060 800
rect 198868 0 198924 800
rect 202640 0 202696 800
rect 206504 0 206560 800
rect 210276 0 210332 800
rect 214048 0 214104 800
rect 217912 0 217968 800
rect 221684 0 221740 800
rect 225548 0 225604 800
rect 229320 0 229376 800
rect 233092 0 233148 800
rect 236956 0 237012 800
rect 240728 0 240784 800
rect 244592 0 244648 800
rect 248364 0 248420 800
rect 252136 0 252192 800
rect 256000 0 256056 800
rect 259772 0 259828 800
rect 263636 0 263692 800
rect 267408 0 267464 800
rect 271180 0 271236 800
rect 275044 0 275100 800
rect 278816 0 278872 800
rect 282680 0 282736 800
rect 286452 0 286508 800
rect 290316 0 290372 800
rect 294088 0 294144 800
rect 297860 0 297916 800
rect 301724 0 301780 800
rect 305496 0 305552 800
rect 309360 0 309416 800
rect 313132 0 313188 800
rect 316904 0 316960 800
rect 320768 0 320824 800
rect 324540 0 324596 800
rect 328404 0 328460 800
rect 332176 0 332232 800
rect 335948 0 336004 800
rect 339812 0 339868 800
rect 343584 0 343640 800
rect 347448 0 347504 800
rect 351220 0 351276 800
rect 354992 0 355048 800
rect 358856 0 358912 800
rect 362628 0 362684 800
rect 366492 0 366548 800
rect 370264 0 370320 800
rect 374128 0 374184 800
rect 377900 0 377956 800
rect 381672 0 381728 800
rect 385536 0 385592 800
rect 389308 0 389364 800
rect 393172 0 393228 800
rect 396944 0 397000 800
rect 400716 0 400772 800
rect 404580 0 404636 800
rect 408352 0 408408 800
rect 412216 0 412272 800
rect 415988 0 416044 800
rect 419760 0 419816 800
rect 423624 0 423680 800
rect 427396 0 427452 800
rect 431260 0 431316 800
rect 435032 0 435088 800
rect 438804 0 438860 800
rect 442668 0 442724 800
rect 446440 0 446496 800
rect 450304 0 450360 800
rect 454076 0 454132 800
rect 457848 0 457904 800
rect 461712 0 461768 800
rect 465484 0 465540 800
rect 469348 0 469404 800
rect 473120 0 473176 800
rect 476984 0 477040 800
rect 480756 0 480812 800
rect 484528 0 484584 800
rect 488392 0 488448 800
rect 492164 0 492220 800
rect 496028 0 496084 800
rect 499800 0 499856 800
rect 503572 0 503628 800
rect 507436 0 507492 800
rect 511208 0 511264 800
rect 515072 0 515128 800
rect 518844 0 518900 800
rect 522616 0 522672 800
rect 526480 0 526536 800
rect 530252 0 530308 800
rect 534116 0 534172 800
rect 537888 0 537944 800
rect 541660 0 541716 800
rect 545524 0 545580 800
rect 549296 0 549352 800
rect 553160 0 553216 800
rect 556932 0 556988 800
<< obsm2 >>
rect 518 856 557354 157808
rect 518 800 736 856
rect 904 800 4508 856
rect 4676 800 8280 856
rect 8448 800 12144 856
rect 12312 800 15916 856
rect 16084 800 19780 856
rect 19948 800 23552 856
rect 23720 800 27324 856
rect 27492 800 31188 856
rect 31356 800 34960 856
rect 35128 800 38824 856
rect 38992 800 42596 856
rect 42764 800 46368 856
rect 46536 800 50232 856
rect 50400 800 54004 856
rect 54172 800 57868 856
rect 58036 800 61640 856
rect 61808 800 65412 856
rect 65580 800 69276 856
rect 69444 800 73048 856
rect 73216 800 76912 856
rect 77080 800 80684 856
rect 80852 800 84456 856
rect 84624 800 88320 856
rect 88488 800 92092 856
rect 92260 800 95956 856
rect 96124 800 99728 856
rect 99896 800 103592 856
rect 103760 800 107364 856
rect 107532 800 111136 856
rect 111304 800 115000 856
rect 115168 800 118772 856
rect 118940 800 122636 856
rect 122804 800 126408 856
rect 126576 800 130180 856
rect 130348 800 134044 856
rect 134212 800 137816 856
rect 137984 800 141680 856
rect 141848 800 145452 856
rect 145620 800 149224 856
rect 149392 800 153088 856
rect 153256 800 156860 856
rect 157028 800 160724 856
rect 160892 800 164496 856
rect 164664 800 168268 856
rect 168436 800 172132 856
rect 172300 800 175904 856
rect 176072 800 179768 856
rect 179936 800 183540 856
rect 183708 800 187404 856
rect 187572 800 191176 856
rect 191344 800 194948 856
rect 195116 800 198812 856
rect 198980 800 202584 856
rect 202752 800 206448 856
rect 206616 800 210220 856
rect 210388 800 213992 856
rect 214160 800 217856 856
rect 218024 800 221628 856
rect 221796 800 225492 856
rect 225660 800 229264 856
rect 229432 800 233036 856
rect 233204 800 236900 856
rect 237068 800 240672 856
rect 240840 800 244536 856
rect 244704 800 248308 856
rect 248476 800 252080 856
rect 252248 800 255944 856
rect 256112 800 259716 856
rect 259884 800 263580 856
rect 263748 800 267352 856
rect 267520 800 271124 856
rect 271292 800 274988 856
rect 275156 800 278760 856
rect 278928 800 282624 856
rect 282792 800 286396 856
rect 286564 800 290260 856
rect 290428 800 294032 856
rect 294200 800 297804 856
rect 297972 800 301668 856
rect 301836 800 305440 856
rect 305608 800 309304 856
rect 309472 800 313076 856
rect 313244 800 316848 856
rect 317016 800 320712 856
rect 320880 800 324484 856
rect 324652 800 328348 856
rect 328516 800 332120 856
rect 332288 800 335892 856
rect 336060 800 339756 856
rect 339924 800 343528 856
rect 343696 800 347392 856
rect 347560 800 351164 856
rect 351332 800 354936 856
rect 355104 800 358800 856
rect 358968 800 362572 856
rect 362740 800 366436 856
rect 366604 800 370208 856
rect 370376 800 374072 856
rect 374240 800 377844 856
rect 378012 800 381616 856
rect 381784 800 385480 856
rect 385648 800 389252 856
rect 389420 800 393116 856
rect 393284 800 396888 856
rect 397056 800 400660 856
rect 400828 800 404524 856
rect 404692 800 408296 856
rect 408464 800 412160 856
rect 412328 800 415932 856
rect 416100 800 419704 856
rect 419872 800 423568 856
rect 423736 800 427340 856
rect 427508 800 431204 856
rect 431372 800 434976 856
rect 435144 800 438748 856
rect 438916 800 442612 856
rect 442780 800 446384 856
rect 446552 800 450248 856
rect 450416 800 454020 856
rect 454188 800 457792 856
rect 457960 800 461656 856
rect 461824 800 465428 856
rect 465596 800 469292 856
rect 469460 800 473064 856
rect 473232 800 476928 856
rect 477096 800 480700 856
rect 480868 800 484472 856
rect 484640 800 488336 856
rect 488504 800 492108 856
rect 492276 800 495972 856
rect 496140 800 499744 856
rect 499912 800 503516 856
rect 503684 800 507380 856
rect 507548 800 511152 856
rect 511320 800 515016 856
rect 515184 800 518788 856
rect 518956 800 522560 856
rect 522728 800 526424 856
rect 526592 800 530196 856
rect 530364 800 534060 856
rect 534228 800 537832 856
rect 538000 800 541604 856
rect 541772 800 545468 856
rect 545636 800 549240 856
rect 549408 800 553104 856
rect 553272 800 556876 856
rect 557044 800 557354 856
<< obsm3 >>
rect 1247 1939 557177 157793
<< metal4 >>
rect 3142 2128 3462 157808
rect 3802 2176 4122 157760
rect 4462 2176 4782 157760
rect 5122 2176 5442 157760
rect 18502 2128 18822 157808
rect 19162 2176 19482 157760
rect 19822 2176 20142 157760
rect 20482 2176 20802 157760
rect 33862 2128 34182 157808
rect 34522 2176 34842 157760
rect 35182 2176 35502 157760
rect 35842 2176 36162 157760
rect 49222 2128 49542 157808
rect 49882 2176 50202 157760
rect 50542 2176 50862 157760
rect 51202 2176 51522 157760
rect 64582 2128 64902 157808
rect 65242 2176 65562 157760
rect 65902 2176 66222 157760
rect 66562 2176 66882 157760
rect 79942 2128 80262 157808
rect 80602 2176 80922 157760
rect 81262 2176 81582 157760
rect 81922 2176 82242 157760
rect 95302 2128 95622 157808
rect 95962 2176 96282 157760
rect 96622 2176 96942 157760
rect 97282 2176 97602 157760
rect 110662 2128 110982 157808
rect 111322 2176 111642 157760
rect 111982 2176 112302 157760
rect 112642 2176 112962 157760
rect 126022 2128 126342 157808
rect 126682 2176 127002 157760
rect 127342 2176 127662 157760
rect 128002 2176 128322 157760
rect 141382 2128 141702 157808
rect 142042 2176 142362 157760
rect 142702 2176 143022 157760
rect 143362 2176 143682 157760
rect 156742 2128 157062 157808
rect 157402 2176 157722 157760
rect 158062 2176 158382 157760
rect 158722 2176 159042 157760
rect 172102 2128 172422 157808
rect 172762 2176 173082 157760
rect 173422 2176 173742 157760
rect 174082 2176 174402 157760
rect 187462 2128 187782 157808
rect 188122 2176 188442 157760
rect 188782 2176 189102 157760
rect 189442 2176 189762 157760
rect 202822 2128 203142 157808
rect 203482 2176 203802 157760
rect 204142 2176 204462 157760
rect 204802 2176 205122 157760
rect 218182 2128 218502 157808
rect 218842 2176 219162 157760
rect 219502 2176 219822 157760
rect 220162 2176 220482 157760
rect 233542 2128 233862 157808
rect 234202 2176 234522 157760
rect 234862 2176 235182 157760
rect 235522 2176 235842 157760
rect 248902 2128 249222 157808
rect 249562 2176 249882 157760
rect 250222 2176 250542 157760
rect 250882 2176 251202 157760
rect 264262 2128 264582 157808
rect 264922 2176 265242 157760
rect 265582 2176 265902 157760
rect 266242 2176 266562 157760
rect 279622 2128 279942 157808
rect 280282 2176 280602 157760
rect 280942 2176 281262 157760
rect 281602 2176 281922 157760
rect 294982 2128 295302 157808
rect 295642 2176 295962 157760
rect 296302 2176 296622 157760
rect 296962 2176 297282 157760
rect 310342 2128 310662 157808
rect 311002 2176 311322 157760
rect 311662 2176 311982 157760
rect 312322 2176 312642 157760
rect 325702 2128 326022 157808
rect 326362 2176 326682 157760
rect 327022 2176 327342 157760
rect 327682 2176 328002 157760
rect 341062 2128 341382 157808
rect 341722 2176 342042 157760
rect 342382 2176 342702 157760
rect 343042 2176 343362 157760
rect 356422 2128 356742 157808
rect 357082 2176 357402 157760
rect 357742 2176 358062 157760
rect 358402 2176 358722 157760
rect 371782 2128 372102 157808
rect 372442 2176 372762 157760
rect 373102 2176 373422 157760
rect 373762 2176 374082 157760
rect 387142 2128 387462 157808
rect 387802 2176 388122 157760
rect 388462 2176 388782 157760
rect 389122 2176 389442 157760
rect 402502 2128 402822 157808
rect 403162 2176 403482 157760
rect 403822 2176 404142 157760
rect 404482 2176 404802 157760
rect 417862 2128 418182 157808
rect 418522 2176 418842 157760
rect 419182 2176 419502 157760
rect 419842 2176 420162 157760
rect 433222 2128 433542 157808
rect 433882 2176 434202 157760
rect 434542 2176 434862 157760
rect 435202 2176 435522 157760
rect 448582 2128 448902 157808
rect 449242 2176 449562 157760
rect 449902 2176 450222 157760
rect 450562 2176 450882 157760
rect 463942 2128 464262 157808
rect 464602 2176 464922 157760
rect 465262 2176 465582 157760
rect 465922 2176 466242 157760
rect 479302 2128 479622 157808
rect 479962 2176 480282 157760
rect 480622 2176 480942 157760
rect 481282 2176 481602 157760
rect 494662 2128 494982 157808
rect 495322 2176 495642 157760
rect 495982 2176 496302 157760
rect 496642 2176 496962 157760
rect 510022 2128 510342 157808
rect 510682 2176 511002 157760
rect 511342 2176 511662 157760
rect 512002 2176 512322 157760
rect 525382 2128 525702 157808
rect 526042 2176 526362 157760
rect 526702 2176 527022 157760
rect 527362 2176 527682 157760
rect 540742 2128 541062 157808
rect 541402 2176 541722 157760
rect 542062 2176 542382 157760
rect 542722 2176 543042 157760
rect 556102 2128 556422 157808
rect 556762 2176 557082 157760
<< obsm4 >>
rect 37449 2048 49142 130253
rect 49622 2096 49802 130253
rect 50282 2096 50462 130253
rect 50942 2096 51122 130253
rect 51602 2096 64502 130253
rect 49622 2048 64502 2096
rect 64982 2096 65162 130253
rect 65642 2096 65822 130253
rect 66302 2096 66482 130253
rect 66962 2096 79862 130253
rect 64982 2048 79862 2096
rect 80342 2096 80522 130253
rect 81002 2096 81182 130253
rect 81662 2096 81842 130253
rect 82322 2096 95222 130253
rect 80342 2048 95222 2096
rect 95702 2096 95882 130253
rect 96362 2096 96542 130253
rect 97022 2096 97202 130253
rect 97682 2096 110582 130253
rect 95702 2048 110582 2096
rect 111062 2096 111242 130253
rect 111722 2096 111902 130253
rect 112382 2096 112562 130253
rect 113042 2096 125942 130253
rect 111062 2048 125942 2096
rect 126422 2096 126602 130253
rect 127082 2096 127262 130253
rect 127742 2096 127922 130253
rect 128402 2096 141302 130253
rect 126422 2048 141302 2096
rect 141782 2096 141962 130253
rect 142442 2096 142622 130253
rect 143102 2096 143282 130253
rect 143762 2096 156662 130253
rect 141782 2048 156662 2096
rect 157142 2096 157322 130253
rect 157802 2096 157982 130253
rect 158462 2096 158642 130253
rect 159122 2096 172022 130253
rect 157142 2048 172022 2096
rect 172502 2096 172682 130253
rect 173162 2096 173342 130253
rect 173822 2096 174002 130253
rect 174482 2096 187382 130253
rect 172502 2048 187382 2096
rect 187862 2096 188042 130253
rect 188522 2096 188702 130253
rect 189182 2096 189362 130253
rect 189842 2096 202742 130253
rect 187862 2048 202742 2096
rect 203222 2096 203402 130253
rect 203882 2096 204062 130253
rect 204542 2096 204722 130253
rect 205202 2096 218102 130253
rect 203222 2048 218102 2096
rect 218582 2096 218762 130253
rect 219242 2096 219422 130253
rect 219902 2096 220082 130253
rect 220562 2096 233462 130253
rect 218582 2048 233462 2096
rect 233942 2096 234122 130253
rect 234602 2096 234782 130253
rect 235262 2096 235442 130253
rect 235922 2096 248822 130253
rect 233942 2048 248822 2096
rect 249302 2096 249482 130253
rect 249962 2096 250142 130253
rect 250622 2096 250802 130253
rect 251282 2096 264182 130253
rect 249302 2048 264182 2096
rect 264662 2096 264842 130253
rect 265322 2096 265502 130253
rect 265982 2096 266162 130253
rect 266642 2096 279542 130253
rect 264662 2048 279542 2096
rect 280022 2096 280202 130253
rect 280682 2096 280862 130253
rect 281342 2096 281522 130253
rect 282002 2096 294902 130253
rect 280022 2048 294902 2096
rect 295382 2096 295562 130253
rect 296042 2096 296222 130253
rect 296702 2096 296882 130253
rect 297362 2096 310262 130253
rect 295382 2048 310262 2096
rect 310742 2096 310922 130253
rect 311402 2096 311582 130253
rect 312062 2096 312242 130253
rect 312722 2096 325622 130253
rect 310742 2048 325622 2096
rect 326102 2096 326282 130253
rect 326762 2096 326942 130253
rect 327422 2096 327602 130253
rect 328082 2096 340982 130253
rect 326102 2048 340982 2096
rect 341462 2096 341642 130253
rect 342122 2096 342302 130253
rect 342782 2096 342962 130253
rect 343442 2096 356342 130253
rect 341462 2048 356342 2096
rect 356822 2096 357002 130253
rect 357482 2096 357662 130253
rect 358142 2096 358322 130253
rect 358802 2096 371702 130253
rect 356822 2048 371702 2096
rect 372182 2096 372362 130253
rect 372842 2096 373022 130253
rect 373502 2096 373682 130253
rect 374162 2096 387062 130253
rect 372182 2048 387062 2096
rect 387542 2096 387722 130253
rect 388202 2096 388382 130253
rect 388862 2096 389042 130253
rect 389522 2096 402422 130253
rect 387542 2048 402422 2096
rect 402902 2096 403082 130253
rect 403562 2096 403742 130253
rect 404222 2096 404402 130253
rect 404882 2096 417782 130253
rect 402902 2048 417782 2096
rect 418262 2096 418442 130253
rect 418922 2096 419102 130253
rect 419582 2096 419762 130253
rect 420242 2096 433142 130253
rect 418262 2048 433142 2096
rect 433622 2096 433802 130253
rect 434282 2096 434462 130253
rect 434942 2096 435122 130253
rect 435602 2096 448502 130253
rect 433622 2048 448502 2096
rect 448982 2096 449162 130253
rect 449642 2096 449822 130253
rect 450302 2096 450482 130253
rect 450962 2096 463862 130253
rect 448982 2048 463862 2096
rect 464342 2096 464522 130253
rect 465002 2096 465182 130253
rect 465662 2096 465842 130253
rect 466322 2096 479222 130253
rect 464342 2048 479222 2096
rect 479702 2096 479882 130253
rect 480362 2096 480542 130253
rect 481022 2096 481202 130253
rect 481682 2096 494582 130253
rect 479702 2048 494582 2096
rect 495062 2096 495242 130253
rect 495722 2096 495902 130253
rect 496382 2096 496562 130253
rect 497042 2096 509942 130253
rect 495062 2048 509942 2096
rect 510422 2096 510602 130253
rect 511082 2096 511262 130253
rect 511742 2096 511922 130253
rect 512402 2096 525302 130253
rect 510422 2048 525302 2096
rect 525782 2096 525962 130253
rect 526442 2096 526622 130253
rect 527102 2096 527282 130253
rect 527762 2096 538547 130253
rect 525782 2048 538547 2096
rect 37449 1939 538547 2048
<< obsm5 >>
rect 278362 19220 451274 83460
<< labels >>
rlabel metal2 s 488392 0 488448 800 6 A[0]
port 1 nsew signal input
rlabel metal2 s 492164 0 492220 800 6 A[1]
port 2 nsew signal input
rlabel metal2 s 496028 0 496084 800 6 A[2]
port 3 nsew signal input
rlabel metal2 s 499800 0 499856 800 6 A[3]
port 4 nsew signal input
rlabel metal2 s 503572 0 503628 800 6 A[4]
port 5 nsew signal input
rlabel metal2 s 507436 0 507492 800 6 A[5]
port 6 nsew signal input
rlabel metal2 s 511208 0 511264 800 6 A[6]
port 7 nsew signal input
rlabel metal2 s 515072 0 515128 800 6 A[7]
port 8 nsew signal input
rlabel metal2 s 518844 0 518900 800 6 A[8]
port 9 nsew signal input
rlabel metal2 s 522616 0 522672 800 6 CLK
port 10 nsew signal input
rlabel metal2 s 244592 0 244648 800 6 Di[0]
port 11 nsew signal input
rlabel metal2 s 282680 0 282736 800 6 Di[10]
port 12 nsew signal input
rlabel metal2 s 286452 0 286508 800 6 Di[11]
port 13 nsew signal input
rlabel metal2 s 290316 0 290372 800 6 Di[12]
port 14 nsew signal input
rlabel metal2 s 294088 0 294144 800 6 Di[13]
port 15 nsew signal input
rlabel metal2 s 297860 0 297916 800 6 Di[14]
port 16 nsew signal input
rlabel metal2 s 301724 0 301780 800 6 Di[15]
port 17 nsew signal input
rlabel metal2 s 305496 0 305552 800 6 Di[16]
port 18 nsew signal input
rlabel metal2 s 309360 0 309416 800 6 Di[17]
port 19 nsew signal input
rlabel metal2 s 313132 0 313188 800 6 Di[18]
port 20 nsew signal input
rlabel metal2 s 316904 0 316960 800 6 Di[19]
port 21 nsew signal input
rlabel metal2 s 248364 0 248420 800 6 Di[1]
port 22 nsew signal input
rlabel metal2 s 320768 0 320824 800 6 Di[20]
port 23 nsew signal input
rlabel metal2 s 324540 0 324596 800 6 Di[21]
port 24 nsew signal input
rlabel metal2 s 328404 0 328460 800 6 Di[22]
port 25 nsew signal input
rlabel metal2 s 332176 0 332232 800 6 Di[23]
port 26 nsew signal input
rlabel metal2 s 335948 0 336004 800 6 Di[24]
port 27 nsew signal input
rlabel metal2 s 339812 0 339868 800 6 Di[25]
port 28 nsew signal input
rlabel metal2 s 343584 0 343640 800 6 Di[26]
port 29 nsew signal input
rlabel metal2 s 347448 0 347504 800 6 Di[27]
port 30 nsew signal input
rlabel metal2 s 351220 0 351276 800 6 Di[28]
port 31 nsew signal input
rlabel metal2 s 354992 0 355048 800 6 Di[29]
port 32 nsew signal input
rlabel metal2 s 252136 0 252192 800 6 Di[2]
port 33 nsew signal input
rlabel metal2 s 358856 0 358912 800 6 Di[30]
port 34 nsew signal input
rlabel metal2 s 362628 0 362684 800 6 Di[31]
port 35 nsew signal input
rlabel metal2 s 366492 0 366548 800 6 Di[32]
port 36 nsew signal input
rlabel metal2 s 370264 0 370320 800 6 Di[33]
port 37 nsew signal input
rlabel metal2 s 374128 0 374184 800 6 Di[34]
port 38 nsew signal input
rlabel metal2 s 377900 0 377956 800 6 Di[35]
port 39 nsew signal input
rlabel metal2 s 381672 0 381728 800 6 Di[36]
port 40 nsew signal input
rlabel metal2 s 385536 0 385592 800 6 Di[37]
port 41 nsew signal input
rlabel metal2 s 389308 0 389364 800 6 Di[38]
port 42 nsew signal input
rlabel metal2 s 393172 0 393228 800 6 Di[39]
port 43 nsew signal input
rlabel metal2 s 256000 0 256056 800 6 Di[3]
port 44 nsew signal input
rlabel metal2 s 396944 0 397000 800 6 Di[40]
port 45 nsew signal input
rlabel metal2 s 400716 0 400772 800 6 Di[41]
port 46 nsew signal input
rlabel metal2 s 404580 0 404636 800 6 Di[42]
port 47 nsew signal input
rlabel metal2 s 408352 0 408408 800 6 Di[43]
port 48 nsew signal input
rlabel metal2 s 412216 0 412272 800 6 Di[44]
port 49 nsew signal input
rlabel metal2 s 415988 0 416044 800 6 Di[45]
port 50 nsew signal input
rlabel metal2 s 419760 0 419816 800 6 Di[46]
port 51 nsew signal input
rlabel metal2 s 423624 0 423680 800 6 Di[47]
port 52 nsew signal input
rlabel metal2 s 427396 0 427452 800 6 Di[48]
port 53 nsew signal input
rlabel metal2 s 431260 0 431316 800 6 Di[49]
port 54 nsew signal input
rlabel metal2 s 259772 0 259828 800 6 Di[4]
port 55 nsew signal input
rlabel metal2 s 435032 0 435088 800 6 Di[50]
port 56 nsew signal input
rlabel metal2 s 438804 0 438860 800 6 Di[51]
port 57 nsew signal input
rlabel metal2 s 442668 0 442724 800 6 Di[52]
port 58 nsew signal input
rlabel metal2 s 446440 0 446496 800 6 Di[53]
port 59 nsew signal input
rlabel metal2 s 450304 0 450360 800 6 Di[54]
port 60 nsew signal input
rlabel metal2 s 454076 0 454132 800 6 Di[55]
port 61 nsew signal input
rlabel metal2 s 457848 0 457904 800 6 Di[56]
port 62 nsew signal input
rlabel metal2 s 461712 0 461768 800 6 Di[57]
port 63 nsew signal input
rlabel metal2 s 465484 0 465540 800 6 Di[58]
port 64 nsew signal input
rlabel metal2 s 469348 0 469404 800 6 Di[59]
port 65 nsew signal input
rlabel metal2 s 263636 0 263692 800 6 Di[5]
port 66 nsew signal input
rlabel metal2 s 473120 0 473176 800 6 Di[60]
port 67 nsew signal input
rlabel metal2 s 476984 0 477040 800 6 Di[61]
port 68 nsew signal input
rlabel metal2 s 480756 0 480812 800 6 Di[62]
port 69 nsew signal input
rlabel metal2 s 484528 0 484584 800 6 Di[63]
port 70 nsew signal input
rlabel metal2 s 267408 0 267464 800 6 Di[6]
port 71 nsew signal input
rlabel metal2 s 271180 0 271236 800 6 Di[7]
port 72 nsew signal input
rlabel metal2 s 275044 0 275100 800 6 Di[8]
port 73 nsew signal input
rlabel metal2 s 278816 0 278872 800 6 Di[9]
port 74 nsew signal input
rlabel metal2 s 792 0 848 800 6 Do[0]
port 75 nsew signal output
rlabel metal2 s 38880 0 38936 800 6 Do[10]
port 76 nsew signal output
rlabel metal2 s 42652 0 42708 800 6 Do[11]
port 77 nsew signal output
rlabel metal2 s 46424 0 46480 800 6 Do[12]
port 78 nsew signal output
rlabel metal2 s 50288 0 50344 800 6 Do[13]
port 79 nsew signal output
rlabel metal2 s 54060 0 54116 800 6 Do[14]
port 80 nsew signal output
rlabel metal2 s 57924 0 57980 800 6 Do[15]
port 81 nsew signal output
rlabel metal2 s 61696 0 61752 800 6 Do[16]
port 82 nsew signal output
rlabel metal2 s 65468 0 65524 800 6 Do[17]
port 83 nsew signal output
rlabel metal2 s 69332 0 69388 800 6 Do[18]
port 84 nsew signal output
rlabel metal2 s 73104 0 73160 800 6 Do[19]
port 85 nsew signal output
rlabel metal2 s 4564 0 4620 800 6 Do[1]
port 86 nsew signal output
rlabel metal2 s 76968 0 77024 800 6 Do[20]
port 87 nsew signal output
rlabel metal2 s 80740 0 80796 800 6 Do[21]
port 88 nsew signal output
rlabel metal2 s 84512 0 84568 800 6 Do[22]
port 89 nsew signal output
rlabel metal2 s 88376 0 88432 800 6 Do[23]
port 90 nsew signal output
rlabel metal2 s 92148 0 92204 800 6 Do[24]
port 91 nsew signal output
rlabel metal2 s 96012 0 96068 800 6 Do[25]
port 92 nsew signal output
rlabel metal2 s 99784 0 99840 800 6 Do[26]
port 93 nsew signal output
rlabel metal2 s 103648 0 103704 800 6 Do[27]
port 94 nsew signal output
rlabel metal2 s 107420 0 107476 800 6 Do[28]
port 95 nsew signal output
rlabel metal2 s 111192 0 111248 800 6 Do[29]
port 96 nsew signal output
rlabel metal2 s 8336 0 8392 800 6 Do[2]
port 97 nsew signal output
rlabel metal2 s 115056 0 115112 800 6 Do[30]
port 98 nsew signal output
rlabel metal2 s 118828 0 118884 800 6 Do[31]
port 99 nsew signal output
rlabel metal2 s 122692 0 122748 800 6 Do[32]
port 100 nsew signal output
rlabel metal2 s 126464 0 126520 800 6 Do[33]
port 101 nsew signal output
rlabel metal2 s 130236 0 130292 800 6 Do[34]
port 102 nsew signal output
rlabel metal2 s 134100 0 134156 800 6 Do[35]
port 103 nsew signal output
rlabel metal2 s 137872 0 137928 800 6 Do[36]
port 104 nsew signal output
rlabel metal2 s 141736 0 141792 800 6 Do[37]
port 105 nsew signal output
rlabel metal2 s 145508 0 145564 800 6 Do[38]
port 106 nsew signal output
rlabel metal2 s 149280 0 149336 800 6 Do[39]
port 107 nsew signal output
rlabel metal2 s 12200 0 12256 800 6 Do[3]
port 108 nsew signal output
rlabel metal2 s 153144 0 153200 800 6 Do[40]
port 109 nsew signal output
rlabel metal2 s 156916 0 156972 800 6 Do[41]
port 110 nsew signal output
rlabel metal2 s 160780 0 160836 800 6 Do[42]
port 111 nsew signal output
rlabel metal2 s 164552 0 164608 800 6 Do[43]
port 112 nsew signal output
rlabel metal2 s 168324 0 168380 800 6 Do[44]
port 113 nsew signal output
rlabel metal2 s 172188 0 172244 800 6 Do[45]
port 114 nsew signal output
rlabel metal2 s 175960 0 176016 800 6 Do[46]
port 115 nsew signal output
rlabel metal2 s 179824 0 179880 800 6 Do[47]
port 116 nsew signal output
rlabel metal2 s 183596 0 183652 800 6 Do[48]
port 117 nsew signal output
rlabel metal2 s 187460 0 187516 800 6 Do[49]
port 118 nsew signal output
rlabel metal2 s 15972 0 16028 800 6 Do[4]
port 119 nsew signal output
rlabel metal2 s 191232 0 191288 800 6 Do[50]
port 120 nsew signal output
rlabel metal2 s 195004 0 195060 800 6 Do[51]
port 121 nsew signal output
rlabel metal2 s 198868 0 198924 800 6 Do[52]
port 122 nsew signal output
rlabel metal2 s 202640 0 202696 800 6 Do[53]
port 123 nsew signal output
rlabel metal2 s 206504 0 206560 800 6 Do[54]
port 124 nsew signal output
rlabel metal2 s 210276 0 210332 800 6 Do[55]
port 125 nsew signal output
rlabel metal2 s 214048 0 214104 800 6 Do[56]
port 126 nsew signal output
rlabel metal2 s 217912 0 217968 800 6 Do[57]
port 127 nsew signal output
rlabel metal2 s 221684 0 221740 800 6 Do[58]
port 128 nsew signal output
rlabel metal2 s 225548 0 225604 800 6 Do[59]
port 129 nsew signal output
rlabel metal2 s 19836 0 19892 800 6 Do[5]
port 130 nsew signal output
rlabel metal2 s 229320 0 229376 800 6 Do[60]
port 131 nsew signal output
rlabel metal2 s 233092 0 233148 800 6 Do[61]
port 132 nsew signal output
rlabel metal2 s 236956 0 237012 800 6 Do[62]
port 133 nsew signal output
rlabel metal2 s 240728 0 240784 800 6 Do[63]
port 134 nsew signal output
rlabel metal2 s 23608 0 23664 800 6 Do[6]
port 135 nsew signal output
rlabel metal2 s 27380 0 27436 800 6 Do[7]
port 136 nsew signal output
rlabel metal2 s 31244 0 31300 800 6 Do[8]
port 137 nsew signal output
rlabel metal2 s 35016 0 35072 800 6 Do[9]
port 138 nsew signal output
rlabel metal2 s 556932 0 556988 800 6 EN
port 139 nsew signal input
rlabel metal2 s 526480 0 526536 800 6 WE[0]
port 140 nsew signal input
rlabel metal2 s 530252 0 530308 800 6 WE[1]
port 141 nsew signal input
rlabel metal2 s 534116 0 534172 800 6 WE[2]
port 142 nsew signal input
rlabel metal2 s 537888 0 537944 800 6 WE[3]
port 143 nsew signal input
rlabel metal2 s 541660 0 541716 800 6 WE[4]
port 144 nsew signal input
rlabel metal2 s 545524 0 545580 800 6 WE[5]
port 145 nsew signal input
rlabel metal2 s 549296 0 549352 800 6 WE[6]
port 146 nsew signal input
rlabel metal2 s 553160 0 553216 800 6 WE[7]
port 147 nsew signal input
rlabel metal4 s 556102 2128 556422 157808 6 vccd1
port 148 nsew power bidirectional
rlabel metal4 s 525382 2128 525702 157808 6 vccd1
port 149 nsew power bidirectional
rlabel metal4 s 494662 2128 494982 157808 6 vccd1
port 150 nsew power bidirectional
rlabel metal4 s 463942 2128 464262 157808 6 vccd1
port 151 nsew power bidirectional
rlabel metal4 s 433222 2128 433542 157808 6 vccd1
port 152 nsew power bidirectional
rlabel metal4 s 402502 2128 402822 157808 6 vccd1
port 153 nsew power bidirectional
rlabel metal4 s 371782 2128 372102 157808 6 vccd1
port 154 nsew power bidirectional
rlabel metal4 s 341062 2128 341382 157808 6 vccd1
port 155 nsew power bidirectional
rlabel metal4 s 310342 2128 310662 157808 6 vccd1
port 156 nsew power bidirectional
rlabel metal4 s 279622 2128 279942 157808 6 vccd1
port 157 nsew power bidirectional
rlabel metal4 s 248902 2128 249222 157808 6 vccd1
port 158 nsew power bidirectional
rlabel metal4 s 218182 2128 218502 157808 6 vccd1
port 159 nsew power bidirectional
rlabel metal4 s 187462 2128 187782 157808 6 vccd1
port 160 nsew power bidirectional
rlabel metal4 s 156742 2128 157062 157808 6 vccd1
port 161 nsew power bidirectional
rlabel metal4 s 126022 2128 126342 157808 6 vccd1
port 162 nsew power bidirectional
rlabel metal4 s 95302 2128 95622 157808 6 vccd1
port 163 nsew power bidirectional
rlabel metal4 s 64582 2128 64902 157808 6 vccd1
port 164 nsew power bidirectional
rlabel metal4 s 33862 2128 34182 157808 6 vccd1
port 165 nsew power bidirectional
rlabel metal4 s 3142 2128 3462 157808 6 vccd1
port 166 nsew power bidirectional
rlabel metal4 s 540742 2128 541062 157808 6 vssd1
port 167 nsew ground bidirectional
rlabel metal4 s 510022 2128 510342 157808 6 vssd1
port 168 nsew ground bidirectional
rlabel metal4 s 479302 2128 479622 157808 6 vssd1
port 169 nsew ground bidirectional
rlabel metal4 s 448582 2128 448902 157808 6 vssd1
port 170 nsew ground bidirectional
rlabel metal4 s 417862 2128 418182 157808 6 vssd1
port 171 nsew ground bidirectional
rlabel metal4 s 387142 2128 387462 157808 6 vssd1
port 172 nsew ground bidirectional
rlabel metal4 s 356422 2128 356742 157808 6 vssd1
port 173 nsew ground bidirectional
rlabel metal4 s 325702 2128 326022 157808 6 vssd1
port 174 nsew ground bidirectional
rlabel metal4 s 294982 2128 295302 157808 6 vssd1
port 175 nsew ground bidirectional
rlabel metal4 s 264262 2128 264582 157808 6 vssd1
port 176 nsew ground bidirectional
rlabel metal4 s 233542 2128 233862 157808 6 vssd1
port 177 nsew ground bidirectional
rlabel metal4 s 202822 2128 203142 157808 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 172102 2128 172422 157808 6 vssd1
port 179 nsew ground bidirectional
rlabel metal4 s 141382 2128 141702 157808 6 vssd1
port 180 nsew ground bidirectional
rlabel metal4 s 110662 2128 110982 157808 6 vssd1
port 181 nsew ground bidirectional
rlabel metal4 s 79942 2128 80262 157808 6 vssd1
port 182 nsew ground bidirectional
rlabel metal4 s 49222 2128 49542 157808 6 vssd1
port 183 nsew ground bidirectional
rlabel metal4 s 18502 2128 18822 157808 6 vssd1
port 184 nsew ground bidirectional
rlabel metal4 s 556762 2176 557082 157760 6 vccd2
port 185 nsew power bidirectional
rlabel metal4 s 526042 2176 526362 157760 6 vccd2
port 186 nsew power bidirectional
rlabel metal4 s 495322 2176 495642 157760 6 vccd2
port 187 nsew power bidirectional
rlabel metal4 s 464602 2176 464922 157760 6 vccd2
port 188 nsew power bidirectional
rlabel metal4 s 433882 2176 434202 157760 6 vccd2
port 189 nsew power bidirectional
rlabel metal4 s 403162 2176 403482 157760 6 vccd2
port 190 nsew power bidirectional
rlabel metal4 s 372442 2176 372762 157760 6 vccd2
port 191 nsew power bidirectional
rlabel metal4 s 341722 2176 342042 157760 6 vccd2
port 192 nsew power bidirectional
rlabel metal4 s 311002 2176 311322 157760 6 vccd2
port 193 nsew power bidirectional
rlabel metal4 s 280282 2176 280602 157760 6 vccd2
port 194 nsew power bidirectional
rlabel metal4 s 249562 2176 249882 157760 6 vccd2
port 195 nsew power bidirectional
rlabel metal4 s 218842 2176 219162 157760 6 vccd2
port 196 nsew power bidirectional
rlabel metal4 s 188122 2176 188442 157760 6 vccd2
port 197 nsew power bidirectional
rlabel metal4 s 157402 2176 157722 157760 6 vccd2
port 198 nsew power bidirectional
rlabel metal4 s 126682 2176 127002 157760 6 vccd2
port 199 nsew power bidirectional
rlabel metal4 s 95962 2176 96282 157760 6 vccd2
port 200 nsew power bidirectional
rlabel metal4 s 65242 2176 65562 157760 6 vccd2
port 201 nsew power bidirectional
rlabel metal4 s 34522 2176 34842 157760 6 vccd2
port 202 nsew power bidirectional
rlabel metal4 s 3802 2176 4122 157760 6 vccd2
port 203 nsew power bidirectional
rlabel metal4 s 541402 2176 541722 157760 6 vssd2
port 204 nsew ground bidirectional
rlabel metal4 s 510682 2176 511002 157760 6 vssd2
port 205 nsew ground bidirectional
rlabel metal4 s 479962 2176 480282 157760 6 vssd2
port 206 nsew ground bidirectional
rlabel metal4 s 449242 2176 449562 157760 6 vssd2
port 207 nsew ground bidirectional
rlabel metal4 s 418522 2176 418842 157760 6 vssd2
port 208 nsew ground bidirectional
rlabel metal4 s 387802 2176 388122 157760 6 vssd2
port 209 nsew ground bidirectional
rlabel metal4 s 357082 2176 357402 157760 6 vssd2
port 210 nsew ground bidirectional
rlabel metal4 s 326362 2176 326682 157760 6 vssd2
port 211 nsew ground bidirectional
rlabel metal4 s 295642 2176 295962 157760 6 vssd2
port 212 nsew ground bidirectional
rlabel metal4 s 264922 2176 265242 157760 6 vssd2
port 213 nsew ground bidirectional
rlabel metal4 s 234202 2176 234522 157760 6 vssd2
port 214 nsew ground bidirectional
rlabel metal4 s 203482 2176 203802 157760 6 vssd2
port 215 nsew ground bidirectional
rlabel metal4 s 172762 2176 173082 157760 6 vssd2
port 216 nsew ground bidirectional
rlabel metal4 s 142042 2176 142362 157760 6 vssd2
port 217 nsew ground bidirectional
rlabel metal4 s 111322 2176 111642 157760 6 vssd2
port 218 nsew ground bidirectional
rlabel metal4 s 80602 2176 80922 157760 6 vssd2
port 219 nsew ground bidirectional
rlabel metal4 s 49882 2176 50202 157760 6 vssd2
port 220 nsew ground bidirectional
rlabel metal4 s 19162 2176 19482 157760 6 vssd2
port 221 nsew ground bidirectional
rlabel metal4 s 526702 2176 527022 157760 6 vdda1
port 222 nsew power bidirectional
rlabel metal4 s 495982 2176 496302 157760 6 vdda1
port 223 nsew power bidirectional
rlabel metal4 s 465262 2176 465582 157760 6 vdda1
port 224 nsew power bidirectional
rlabel metal4 s 434542 2176 434862 157760 6 vdda1
port 225 nsew power bidirectional
rlabel metal4 s 403822 2176 404142 157760 6 vdda1
port 226 nsew power bidirectional
rlabel metal4 s 373102 2176 373422 157760 6 vdda1
port 227 nsew power bidirectional
rlabel metal4 s 342382 2176 342702 157760 6 vdda1
port 228 nsew power bidirectional
rlabel metal4 s 311662 2176 311982 157760 6 vdda1
port 229 nsew power bidirectional
rlabel metal4 s 280942 2176 281262 157760 6 vdda1
port 230 nsew power bidirectional
rlabel metal4 s 250222 2176 250542 157760 6 vdda1
port 231 nsew power bidirectional
rlabel metal4 s 219502 2176 219822 157760 6 vdda1
port 232 nsew power bidirectional
rlabel metal4 s 188782 2176 189102 157760 6 vdda1
port 233 nsew power bidirectional
rlabel metal4 s 158062 2176 158382 157760 6 vdda1
port 234 nsew power bidirectional
rlabel metal4 s 127342 2176 127662 157760 6 vdda1
port 235 nsew power bidirectional
rlabel metal4 s 96622 2176 96942 157760 6 vdda1
port 236 nsew power bidirectional
rlabel metal4 s 65902 2176 66222 157760 6 vdda1
port 237 nsew power bidirectional
rlabel metal4 s 35182 2176 35502 157760 6 vdda1
port 238 nsew power bidirectional
rlabel metal4 s 4462 2176 4782 157760 6 vdda1
port 239 nsew power bidirectional
rlabel metal4 s 542062 2176 542382 157760 6 vssa1
port 240 nsew ground bidirectional
rlabel metal4 s 511342 2176 511662 157760 6 vssa1
port 241 nsew ground bidirectional
rlabel metal4 s 480622 2176 480942 157760 6 vssa1
port 242 nsew ground bidirectional
rlabel metal4 s 449902 2176 450222 157760 6 vssa1
port 243 nsew ground bidirectional
rlabel metal4 s 419182 2176 419502 157760 6 vssa1
port 244 nsew ground bidirectional
rlabel metal4 s 388462 2176 388782 157760 6 vssa1
port 245 nsew ground bidirectional
rlabel metal4 s 357742 2176 358062 157760 6 vssa1
port 246 nsew ground bidirectional
rlabel metal4 s 327022 2176 327342 157760 6 vssa1
port 247 nsew ground bidirectional
rlabel metal4 s 296302 2176 296622 157760 6 vssa1
port 248 nsew ground bidirectional
rlabel metal4 s 265582 2176 265902 157760 6 vssa1
port 249 nsew ground bidirectional
rlabel metal4 s 234862 2176 235182 157760 6 vssa1
port 250 nsew ground bidirectional
rlabel metal4 s 204142 2176 204462 157760 6 vssa1
port 251 nsew ground bidirectional
rlabel metal4 s 173422 2176 173742 157760 6 vssa1
port 252 nsew ground bidirectional
rlabel metal4 s 142702 2176 143022 157760 6 vssa1
port 253 nsew ground bidirectional
rlabel metal4 s 111982 2176 112302 157760 6 vssa1
port 254 nsew ground bidirectional
rlabel metal4 s 81262 2176 81582 157760 6 vssa1
port 255 nsew ground bidirectional
rlabel metal4 s 50542 2176 50862 157760 6 vssa1
port 256 nsew ground bidirectional
rlabel metal4 s 19822 2176 20142 157760 6 vssa1
port 257 nsew ground bidirectional
rlabel metal4 s 527362 2176 527682 157760 6 vdda2
port 258 nsew power bidirectional
rlabel metal4 s 496642 2176 496962 157760 6 vdda2
port 259 nsew power bidirectional
rlabel metal4 s 465922 2176 466242 157760 6 vdda2
port 260 nsew power bidirectional
rlabel metal4 s 435202 2176 435522 157760 6 vdda2
port 261 nsew power bidirectional
rlabel metal4 s 404482 2176 404802 157760 6 vdda2
port 262 nsew power bidirectional
rlabel metal4 s 373762 2176 374082 157760 6 vdda2
port 263 nsew power bidirectional
rlabel metal4 s 343042 2176 343362 157760 6 vdda2
port 264 nsew power bidirectional
rlabel metal4 s 312322 2176 312642 157760 6 vdda2
port 265 nsew power bidirectional
rlabel metal4 s 281602 2176 281922 157760 6 vdda2
port 266 nsew power bidirectional
rlabel metal4 s 250882 2176 251202 157760 6 vdda2
port 267 nsew power bidirectional
rlabel metal4 s 220162 2176 220482 157760 6 vdda2
port 268 nsew power bidirectional
rlabel metal4 s 189442 2176 189762 157760 6 vdda2
port 269 nsew power bidirectional
rlabel metal4 s 158722 2176 159042 157760 6 vdda2
port 270 nsew power bidirectional
rlabel metal4 s 128002 2176 128322 157760 6 vdda2
port 271 nsew power bidirectional
rlabel metal4 s 97282 2176 97602 157760 6 vdda2
port 272 nsew power bidirectional
rlabel metal4 s 66562 2176 66882 157760 6 vdda2
port 273 nsew power bidirectional
rlabel metal4 s 35842 2176 36162 157760 6 vdda2
port 274 nsew power bidirectional
rlabel metal4 s 5122 2176 5442 157760 6 vdda2
port 275 nsew power bidirectional
rlabel metal4 s 542722 2176 543042 157760 6 vssa2
port 276 nsew ground bidirectional
rlabel metal4 s 512002 2176 512322 157760 6 vssa2
port 277 nsew ground bidirectional
rlabel metal4 s 481282 2176 481602 157760 6 vssa2
port 278 nsew ground bidirectional
rlabel metal4 s 450562 2176 450882 157760 6 vssa2
port 279 nsew ground bidirectional
rlabel metal4 s 419842 2176 420162 157760 6 vssa2
port 280 nsew ground bidirectional
rlabel metal4 s 389122 2176 389442 157760 6 vssa2
port 281 nsew ground bidirectional
rlabel metal4 s 358402 2176 358722 157760 6 vssa2
port 282 nsew ground bidirectional
rlabel metal4 s 327682 2176 328002 157760 6 vssa2
port 283 nsew ground bidirectional
rlabel metal4 s 296962 2176 297282 157760 6 vssa2
port 284 nsew ground bidirectional
rlabel metal4 s 266242 2176 266562 157760 6 vssa2
port 285 nsew ground bidirectional
rlabel metal4 s 235522 2176 235842 157760 6 vssa2
port 286 nsew ground bidirectional
rlabel metal4 s 204802 2176 205122 157760 6 vssa2
port 287 nsew ground bidirectional
rlabel metal4 s 174082 2176 174402 157760 6 vssa2
port 288 nsew ground bidirectional
rlabel metal4 s 143362 2176 143682 157760 6 vssa2
port 289 nsew ground bidirectional
rlabel metal4 s 112642 2176 112962 157760 6 vssa2
port 290 nsew ground bidirectional
rlabel metal4 s 81922 2176 82242 157760 6 vssa2
port 291 nsew ground bidirectional
rlabel metal4 s 51202 2176 51522 157760 6 vssa2
port 292 nsew ground bidirectional
rlabel metal4 s 20482 2176 20802 157760 6 vssa2
port 293 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 557780 157808
string LEFview TRUE
<< end >>
