magic
tech sky130A
magscale 1 2
timestamp 1608837633
<< obsli1 >>
rect 722 1377 130442 129489
<< obsm1 >>
rect 0 8 131256 131164
<< metal2 >>
rect 4 131200 60 132000
rect 740 131200 796 132000
rect 1476 131200 1532 132000
rect 2212 131200 2268 132000
rect 3040 131200 3096 132000
rect 3776 131200 3832 132000
rect 4512 131200 4568 132000
rect 5340 131200 5396 132000
rect 6076 131200 6132 132000
rect 6812 131200 6868 132000
rect 7548 131200 7604 132000
rect 8376 131200 8432 132000
rect 9112 131200 9168 132000
rect 9848 131200 9904 132000
rect 10676 131200 10732 132000
rect 11412 131200 11468 132000
rect 12148 131200 12204 132000
rect 12976 131200 13032 132000
rect 13712 131200 13768 132000
rect 14448 131200 14504 132000
rect 15184 131200 15240 132000
rect 16012 131200 16068 132000
rect 16748 131200 16804 132000
rect 17484 131200 17540 132000
rect 18312 131200 18368 132000
rect 19048 131200 19104 132000
rect 19784 131200 19840 132000
rect 20520 131200 20576 132000
rect 21348 131200 21404 132000
rect 22084 131200 22140 132000
rect 22820 131200 22876 132000
rect 23648 131200 23704 132000
rect 24384 131200 24440 132000
rect 25120 131200 25176 132000
rect 25948 131200 26004 132000
rect 26684 131200 26740 132000
rect 27420 131200 27476 132000
rect 28156 131200 28212 132000
rect 28984 131200 29040 132000
rect 29720 131200 29776 132000
rect 30456 131200 30512 132000
rect 31284 131200 31340 132000
rect 32020 131200 32076 132000
rect 32756 131200 32812 132000
rect 33492 131200 33548 132000
rect 34320 131200 34376 132000
rect 35056 131200 35112 132000
rect 35792 131200 35848 132000
rect 36620 131200 36676 132000
rect 37356 131200 37412 132000
rect 38092 131200 38148 132000
rect 38920 131200 38976 132000
rect 39656 131200 39712 132000
rect 40392 131200 40448 132000
rect 41128 131200 41184 132000
rect 41956 131200 42012 132000
rect 42692 131200 42748 132000
rect 43428 131200 43484 132000
rect 44256 131200 44312 132000
rect 44992 131200 45048 132000
rect 45728 131200 45784 132000
rect 46464 131200 46520 132000
rect 47292 131200 47348 132000
rect 48028 131200 48084 132000
rect 48764 131200 48820 132000
rect 49592 131200 49648 132000
rect 50328 131200 50384 132000
rect 51064 131200 51120 132000
rect 51892 131200 51948 132000
rect 52628 131200 52684 132000
rect 53364 131200 53420 132000
rect 54100 131200 54156 132000
rect 54928 131200 54984 132000
rect 55664 131200 55720 132000
rect 56400 131200 56456 132000
rect 57228 131200 57284 132000
rect 57964 131200 58020 132000
rect 58700 131200 58756 132000
rect 59436 131200 59492 132000
rect 60264 131200 60320 132000
rect 61000 131200 61056 132000
rect 61736 131200 61792 132000
rect 62564 131200 62620 132000
rect 63300 131200 63356 132000
rect 64036 131200 64092 132000
rect 64864 131200 64920 132000
rect 65600 131200 65656 132000
rect 66336 131200 66392 132000
rect 67072 131200 67128 132000
rect 67900 131200 67956 132000
rect 68636 131200 68692 132000
rect 69372 131200 69428 132000
rect 70200 131200 70256 132000
rect 70936 131200 70992 132000
rect 71672 131200 71728 132000
rect 72500 131200 72556 132000
rect 73236 131200 73292 132000
rect 73972 131200 74028 132000
rect 74708 131200 74764 132000
rect 75536 131200 75592 132000
rect 76272 131200 76328 132000
rect 77008 131200 77064 132000
rect 77836 131200 77892 132000
rect 78572 131200 78628 132000
rect 79308 131200 79364 132000
rect 80044 131200 80100 132000
rect 80872 131200 80928 132000
rect 81608 131200 81664 132000
rect 82344 131200 82400 132000
rect 83172 131200 83228 132000
rect 83908 131200 83964 132000
rect 84644 131200 84700 132000
rect 85472 131200 85528 132000
rect 86208 131200 86264 132000
rect 86944 131200 87000 132000
rect 87680 131200 87736 132000
rect 88508 131200 88564 132000
rect 89244 131200 89300 132000
rect 89980 131200 90036 132000
rect 90808 131200 90864 132000
rect 91544 131200 91600 132000
rect 92280 131200 92336 132000
rect 93016 131200 93072 132000
rect 93844 131200 93900 132000
rect 94580 131200 94636 132000
rect 95316 131200 95372 132000
rect 96144 131200 96200 132000
rect 96880 131200 96936 132000
rect 97616 131200 97672 132000
rect 98444 131200 98500 132000
rect 99180 131200 99236 132000
rect 99916 131200 99972 132000
rect 100652 131200 100708 132000
rect 101480 131200 101536 132000
rect 102216 131200 102272 132000
rect 102952 131200 103008 132000
rect 103780 131200 103836 132000
rect 104516 131200 104572 132000
rect 105252 131200 105308 132000
rect 105988 131200 106044 132000
rect 106816 131200 106872 132000
rect 107552 131200 107608 132000
rect 108288 131200 108344 132000
rect 109116 131200 109172 132000
rect 109852 131200 109908 132000
rect 110588 131200 110644 132000
rect 111416 131200 111472 132000
rect 112152 131200 112208 132000
rect 112888 131200 112944 132000
rect 113624 131200 113680 132000
rect 114452 131200 114508 132000
rect 115188 131200 115244 132000
rect 115924 131200 115980 132000
rect 116752 131200 116808 132000
rect 117488 131200 117544 132000
rect 118224 131200 118280 132000
rect 118960 131200 119016 132000
rect 119788 131200 119844 132000
rect 120524 131200 120580 132000
rect 121260 131200 121316 132000
rect 122088 131200 122144 132000
rect 122824 131200 122880 132000
rect 123560 131200 123616 132000
rect 124388 131200 124444 132000
rect 125124 131200 125180 132000
rect 125860 131200 125916 132000
rect 126596 131200 126652 132000
rect 127424 131200 127480 132000
rect 128160 131200 128216 132000
rect 128896 131200 128952 132000
rect 129724 131200 129780 132000
rect 130460 131200 130516 132000
rect 131196 131200 131252 132000
rect 4 0 60 800
rect 740 0 796 800
rect 1476 0 1532 800
rect 2212 0 2268 800
rect 3040 0 3096 800
rect 3776 0 3832 800
rect 4512 0 4568 800
rect 5340 0 5396 800
rect 6076 0 6132 800
rect 6812 0 6868 800
rect 7548 0 7604 800
rect 8376 0 8432 800
rect 9112 0 9168 800
rect 9848 0 9904 800
rect 10676 0 10732 800
rect 11412 0 11468 800
rect 12148 0 12204 800
rect 12976 0 13032 800
rect 13712 0 13768 800
rect 14448 0 14504 800
rect 15184 0 15240 800
rect 16012 0 16068 800
rect 16748 0 16804 800
rect 17484 0 17540 800
rect 18312 0 18368 800
rect 19048 0 19104 800
rect 19784 0 19840 800
rect 20520 0 20576 800
rect 21348 0 21404 800
rect 22084 0 22140 800
rect 22820 0 22876 800
rect 23648 0 23704 800
rect 24384 0 24440 800
rect 25120 0 25176 800
rect 25948 0 26004 800
rect 26684 0 26740 800
rect 27420 0 27476 800
rect 28156 0 28212 800
rect 28984 0 29040 800
rect 29720 0 29776 800
rect 30456 0 30512 800
rect 31284 0 31340 800
rect 32020 0 32076 800
rect 32756 0 32812 800
rect 33492 0 33548 800
rect 34320 0 34376 800
rect 35056 0 35112 800
rect 35792 0 35848 800
rect 36620 0 36676 800
rect 37356 0 37412 800
rect 38092 0 38148 800
rect 38920 0 38976 800
rect 39656 0 39712 800
rect 40392 0 40448 800
rect 41128 0 41184 800
rect 41956 0 42012 800
rect 42692 0 42748 800
rect 43428 0 43484 800
rect 44256 0 44312 800
rect 44992 0 45048 800
rect 45728 0 45784 800
rect 46464 0 46520 800
rect 47292 0 47348 800
rect 48028 0 48084 800
rect 48764 0 48820 800
rect 49592 0 49648 800
rect 50328 0 50384 800
rect 51064 0 51120 800
rect 51892 0 51948 800
rect 52628 0 52684 800
rect 53364 0 53420 800
rect 54100 0 54156 800
rect 54928 0 54984 800
rect 55664 0 55720 800
rect 56400 0 56456 800
rect 57228 0 57284 800
rect 57964 0 58020 800
rect 58700 0 58756 800
rect 59436 0 59492 800
rect 60264 0 60320 800
rect 61000 0 61056 800
rect 61736 0 61792 800
rect 62564 0 62620 800
rect 63300 0 63356 800
rect 64036 0 64092 800
rect 64864 0 64920 800
rect 65600 0 65656 800
rect 66336 0 66392 800
rect 67072 0 67128 800
rect 67900 0 67956 800
rect 68636 0 68692 800
rect 69372 0 69428 800
rect 70200 0 70256 800
rect 70936 0 70992 800
rect 71672 0 71728 800
rect 72500 0 72556 800
rect 73236 0 73292 800
rect 73972 0 74028 800
rect 74708 0 74764 800
rect 75536 0 75592 800
rect 76272 0 76328 800
rect 77008 0 77064 800
rect 77836 0 77892 800
rect 78572 0 78628 800
rect 79308 0 79364 800
rect 80044 0 80100 800
rect 80872 0 80928 800
rect 81608 0 81664 800
rect 82344 0 82400 800
rect 83172 0 83228 800
rect 83908 0 83964 800
rect 84644 0 84700 800
rect 85472 0 85528 800
rect 86208 0 86264 800
rect 86944 0 87000 800
rect 87680 0 87736 800
rect 88508 0 88564 800
rect 89244 0 89300 800
rect 89980 0 90036 800
rect 90808 0 90864 800
rect 91544 0 91600 800
rect 92280 0 92336 800
rect 93016 0 93072 800
rect 93844 0 93900 800
rect 94580 0 94636 800
rect 95316 0 95372 800
rect 96144 0 96200 800
rect 96880 0 96936 800
rect 97616 0 97672 800
rect 98444 0 98500 800
rect 99180 0 99236 800
rect 99916 0 99972 800
rect 100652 0 100708 800
rect 101480 0 101536 800
rect 102216 0 102272 800
rect 102952 0 103008 800
rect 103780 0 103836 800
rect 104516 0 104572 800
rect 105252 0 105308 800
rect 105988 0 106044 800
rect 106816 0 106872 800
rect 107552 0 107608 800
rect 108288 0 108344 800
rect 109116 0 109172 800
rect 109852 0 109908 800
rect 110588 0 110644 800
rect 111416 0 111472 800
rect 112152 0 112208 800
rect 112888 0 112944 800
rect 113624 0 113680 800
rect 114452 0 114508 800
rect 115188 0 115244 800
rect 115924 0 115980 800
rect 116752 0 116808 800
rect 117488 0 117544 800
rect 118224 0 118280 800
rect 118960 0 119016 800
rect 119788 0 119844 800
rect 120524 0 120580 800
rect 121260 0 121316 800
rect 122088 0 122144 800
rect 122824 0 122880 800
rect 123560 0 123616 800
rect 124388 0 124444 800
rect 125124 0 125180 800
rect 125860 0 125916 800
rect 126596 0 126652 800
rect 127424 0 127480 800
rect 128160 0 128216 800
rect 128896 0 128952 800
rect 129724 0 129780 800
rect 130460 0 130516 800
rect 131196 0 131252 800
<< obsm2 >>
rect 116 131144 684 131200
rect 852 131144 1420 131200
rect 1588 131144 2156 131200
rect 2324 131144 2984 131200
rect 3152 131144 3720 131200
rect 3888 131144 4456 131200
rect 4624 131144 5284 131200
rect 5452 131144 6020 131200
rect 6188 131144 6756 131200
rect 6924 131144 7492 131200
rect 7660 131144 8320 131200
rect 8488 131144 9056 131200
rect 9224 131144 9792 131200
rect 9960 131144 10620 131200
rect 10788 131144 11356 131200
rect 11524 131144 12092 131200
rect 12260 131144 12920 131200
rect 13088 131144 13656 131200
rect 13824 131144 14392 131200
rect 14560 131144 15128 131200
rect 15296 131144 15956 131200
rect 16124 131144 16692 131200
rect 16860 131144 17428 131200
rect 17596 131144 18256 131200
rect 18424 131144 18992 131200
rect 19160 131144 19728 131200
rect 19896 131144 20464 131200
rect 20632 131144 21292 131200
rect 21460 131144 22028 131200
rect 22196 131144 22764 131200
rect 22932 131144 23592 131200
rect 23760 131144 24328 131200
rect 24496 131144 25064 131200
rect 25232 131144 25892 131200
rect 26060 131144 26628 131200
rect 26796 131144 27364 131200
rect 27532 131144 28100 131200
rect 28268 131144 28928 131200
rect 29096 131144 29664 131200
rect 29832 131144 30400 131200
rect 30568 131144 31228 131200
rect 31396 131144 31964 131200
rect 32132 131144 32700 131200
rect 32868 131144 33436 131200
rect 33604 131144 34264 131200
rect 34432 131144 35000 131200
rect 35168 131144 35736 131200
rect 35904 131144 36564 131200
rect 36732 131144 37300 131200
rect 37468 131144 38036 131200
rect 38204 131144 38864 131200
rect 39032 131144 39600 131200
rect 39768 131144 40336 131200
rect 40504 131144 41072 131200
rect 41240 131144 41900 131200
rect 42068 131144 42636 131200
rect 42804 131144 43372 131200
rect 43540 131144 44200 131200
rect 44368 131144 44936 131200
rect 45104 131144 45672 131200
rect 45840 131144 46408 131200
rect 46576 131144 47236 131200
rect 47404 131144 47972 131200
rect 48140 131144 48708 131200
rect 48876 131144 49536 131200
rect 49704 131144 50272 131200
rect 50440 131144 51008 131200
rect 51176 131144 51836 131200
rect 52004 131144 52572 131200
rect 52740 131144 53308 131200
rect 53476 131144 54044 131200
rect 54212 131144 54872 131200
rect 55040 131144 55608 131200
rect 55776 131144 56344 131200
rect 56512 131144 57172 131200
rect 57340 131144 57908 131200
rect 58076 131144 58644 131200
rect 58812 131144 59380 131200
rect 59548 131144 60208 131200
rect 60376 131144 60944 131200
rect 61112 131144 61680 131200
rect 61848 131144 62508 131200
rect 62676 131144 63244 131200
rect 63412 131144 63980 131200
rect 64148 131144 64808 131200
rect 64976 131144 65544 131200
rect 65712 131144 66280 131200
rect 66448 131144 67016 131200
rect 67184 131144 67844 131200
rect 68012 131144 68580 131200
rect 68748 131144 69316 131200
rect 69484 131144 70144 131200
rect 70312 131144 70880 131200
rect 71048 131144 71616 131200
rect 71784 131144 72444 131200
rect 72612 131144 73180 131200
rect 73348 131144 73916 131200
rect 74084 131144 74652 131200
rect 74820 131144 75480 131200
rect 75648 131144 76216 131200
rect 76384 131144 76952 131200
rect 77120 131144 77780 131200
rect 77948 131144 78516 131200
rect 78684 131144 79252 131200
rect 79420 131144 79988 131200
rect 80156 131144 80816 131200
rect 80984 131144 81552 131200
rect 81720 131144 82288 131200
rect 82456 131144 83116 131200
rect 83284 131144 83852 131200
rect 84020 131144 84588 131200
rect 84756 131144 85416 131200
rect 85584 131144 86152 131200
rect 86320 131144 86888 131200
rect 87056 131144 87624 131200
rect 87792 131144 88452 131200
rect 88620 131144 89188 131200
rect 89356 131144 89924 131200
rect 90092 131144 90752 131200
rect 90920 131144 91488 131200
rect 91656 131144 92224 131200
rect 92392 131144 92960 131200
rect 93128 131144 93788 131200
rect 93956 131144 94524 131200
rect 94692 131144 95260 131200
rect 95428 131144 96088 131200
rect 96256 131144 96824 131200
rect 96992 131144 97560 131200
rect 97728 131144 98388 131200
rect 98556 131144 99124 131200
rect 99292 131144 99860 131200
rect 100028 131144 100596 131200
rect 100764 131144 101424 131200
rect 101592 131144 102160 131200
rect 102328 131144 102896 131200
rect 103064 131144 103724 131200
rect 103892 131144 104460 131200
rect 104628 131144 105196 131200
rect 105364 131144 105932 131200
rect 106100 131144 106760 131200
rect 106928 131144 107496 131200
rect 107664 131144 108232 131200
rect 108400 131144 109060 131200
rect 109228 131144 109796 131200
rect 109964 131144 110532 131200
rect 110700 131144 111360 131200
rect 111528 131144 112096 131200
rect 112264 131144 112832 131200
rect 113000 131144 113568 131200
rect 113736 131144 114396 131200
rect 114564 131144 115132 131200
rect 115300 131144 115868 131200
rect 116036 131144 116696 131200
rect 116864 131144 117432 131200
rect 117600 131144 118168 131200
rect 118336 131144 118904 131200
rect 119072 131144 119732 131200
rect 119900 131144 120468 131200
rect 120636 131144 121204 131200
rect 121372 131144 122032 131200
rect 122200 131144 122768 131200
rect 122936 131144 123504 131200
rect 123672 131144 124332 131200
rect 124500 131144 125068 131200
rect 125236 131144 125804 131200
rect 125972 131144 126540 131200
rect 126708 131144 127368 131200
rect 127536 131144 128104 131200
rect 128272 131144 128840 131200
rect 129008 131144 129668 131200
rect 129836 131144 130404 131200
rect 130572 131144 131140 131200
rect 6 856 131250 131144
rect 116 2 684 856
rect 852 2 1420 856
rect 1588 2 2156 856
rect 2324 2 2984 856
rect 3152 2 3720 856
rect 3888 2 4456 856
rect 4624 2 5284 856
rect 5452 2 6020 856
rect 6188 2 6756 856
rect 6924 2 7492 856
rect 7660 2 8320 856
rect 8488 2 9056 856
rect 9224 2 9792 856
rect 9960 2 10620 856
rect 10788 2 11356 856
rect 11524 2 12092 856
rect 12260 2 12920 856
rect 13088 2 13656 856
rect 13824 2 14392 856
rect 14560 2 15128 856
rect 15296 2 15956 856
rect 16124 2 16692 856
rect 16860 2 17428 856
rect 17596 2 18256 856
rect 18424 2 18992 856
rect 19160 2 19728 856
rect 19896 2 20464 856
rect 20632 2 21292 856
rect 21460 2 22028 856
rect 22196 2 22764 856
rect 22932 2 23592 856
rect 23760 2 24328 856
rect 24496 2 25064 856
rect 25232 2 25892 856
rect 26060 2 26628 856
rect 26796 2 27364 856
rect 27532 2 28100 856
rect 28268 2 28928 856
rect 29096 2 29664 856
rect 29832 2 30400 856
rect 30568 2 31228 856
rect 31396 2 31964 856
rect 32132 2 32700 856
rect 32868 2 33436 856
rect 33604 2 34264 856
rect 34432 2 35000 856
rect 35168 2 35736 856
rect 35904 2 36564 856
rect 36732 2 37300 856
rect 37468 2 38036 856
rect 38204 2 38864 856
rect 39032 2 39600 856
rect 39768 2 40336 856
rect 40504 2 41072 856
rect 41240 2 41900 856
rect 42068 2 42636 856
rect 42804 2 43372 856
rect 43540 2 44200 856
rect 44368 2 44936 856
rect 45104 2 45672 856
rect 45840 2 46408 856
rect 46576 2 47236 856
rect 47404 2 47972 856
rect 48140 2 48708 856
rect 48876 2 49536 856
rect 49704 2 50272 856
rect 50440 2 51008 856
rect 51176 2 51836 856
rect 52004 2 52572 856
rect 52740 2 53308 856
rect 53476 2 54044 856
rect 54212 2 54872 856
rect 55040 2 55608 856
rect 55776 2 56344 856
rect 56512 2 57172 856
rect 57340 2 57908 856
rect 58076 2 58644 856
rect 58812 2 59380 856
rect 59548 2 60208 856
rect 60376 2 60944 856
rect 61112 2 61680 856
rect 61848 2 62508 856
rect 62676 2 63244 856
rect 63412 2 63980 856
rect 64148 2 64808 856
rect 64976 2 65544 856
rect 65712 2 66280 856
rect 66448 2 67016 856
rect 67184 2 67844 856
rect 68012 2 68580 856
rect 68748 2 69316 856
rect 69484 2 70144 856
rect 70312 2 70880 856
rect 71048 2 71616 856
rect 71784 2 72444 856
rect 72612 2 73180 856
rect 73348 2 73916 856
rect 74084 2 74652 856
rect 74820 2 75480 856
rect 75648 2 76216 856
rect 76384 2 76952 856
rect 77120 2 77780 856
rect 77948 2 78516 856
rect 78684 2 79252 856
rect 79420 2 79988 856
rect 80156 2 80816 856
rect 80984 2 81552 856
rect 81720 2 82288 856
rect 82456 2 83116 856
rect 83284 2 83852 856
rect 84020 2 84588 856
rect 84756 2 85416 856
rect 85584 2 86152 856
rect 86320 2 86888 856
rect 87056 2 87624 856
rect 87792 2 88452 856
rect 88620 2 89188 856
rect 89356 2 89924 856
rect 90092 2 90752 856
rect 90920 2 91488 856
rect 91656 2 92224 856
rect 92392 2 92960 856
rect 93128 2 93788 856
rect 93956 2 94524 856
rect 94692 2 95260 856
rect 95428 2 96088 856
rect 96256 2 96824 856
rect 96992 2 97560 856
rect 97728 2 98388 856
rect 98556 2 99124 856
rect 99292 2 99860 856
rect 100028 2 100596 856
rect 100764 2 101424 856
rect 101592 2 102160 856
rect 102328 2 102896 856
rect 103064 2 103724 856
rect 103892 2 104460 856
rect 104628 2 105196 856
rect 105364 2 105932 856
rect 106100 2 106760 856
rect 106928 2 107496 856
rect 107664 2 108232 856
rect 108400 2 109060 856
rect 109228 2 109796 856
rect 109964 2 110532 856
rect 110700 2 111360 856
rect 111528 2 112096 856
rect 112264 2 112832 856
rect 113000 2 113568 856
rect 113736 2 114396 856
rect 114564 2 115132 856
rect 115300 2 115868 856
rect 116036 2 116696 856
rect 116864 2 117432 856
rect 117600 2 118168 856
rect 118336 2 118904 856
rect 119072 2 119732 856
rect 119900 2 120468 856
rect 120636 2 121204 856
rect 121372 2 122032 856
rect 122200 2 122768 856
rect 122936 2 123504 856
rect 123672 2 124332 856
rect 124500 2 125068 856
rect 125236 2 125804 856
rect 125972 2 126540 856
rect 126708 2 127368 856
rect 127536 2 128104 856
rect 128272 2 128840 856
rect 129008 2 129668 856
rect 129836 2 130404 856
rect 130572 2 131140 856
<< metal3 >>
rect 130818 131384 131618 131504
rect 130818 130432 131618 130552
rect 130818 129480 131618 129600
rect 130818 128392 131618 128512
rect 130818 127440 131618 127560
rect 130818 126488 131618 126608
rect 130818 125400 131618 125520
rect 130818 124448 131618 124568
rect 130818 123496 131618 123616
rect 130818 122408 131618 122528
rect 130818 121456 131618 121576
rect 130818 120504 131618 120624
rect 130818 119552 131618 119672
rect 130818 118464 131618 118584
rect 130818 117512 131618 117632
rect 130818 116560 131618 116680
rect 130818 115472 131618 115592
rect 130818 114520 131618 114640
rect 130818 113568 131618 113688
rect 130818 112480 131618 112600
rect 130818 111528 131618 111648
rect 130818 110576 131618 110696
rect 130818 109624 131618 109744
rect 130818 108536 131618 108656
rect 130818 107584 131618 107704
rect 130818 106632 131618 106752
rect 130818 105544 131618 105664
rect 130818 104592 131618 104712
rect 130818 103640 131618 103760
rect 130818 102552 131618 102672
rect 130818 101600 131618 101720
rect 130818 100648 131618 100768
rect 130818 99696 131618 99816
rect 130818 98608 131618 98728
rect 130818 97656 131618 97776
rect 130818 96704 131618 96824
rect 130818 95616 131618 95736
rect 130818 94664 131618 94784
rect 130818 93712 131618 93832
rect 130818 92624 131618 92744
rect 130818 91672 131618 91792
rect 130818 90720 131618 90840
rect 130818 89768 131618 89888
rect 130818 88680 131618 88800
rect 130818 87728 131618 87848
rect 130818 86776 131618 86896
rect 130818 85688 131618 85808
rect 130818 84736 131618 84856
rect 130818 83784 131618 83904
rect 130818 82696 131618 82816
rect 130818 81744 131618 81864
rect 130818 80792 131618 80912
rect 130818 79840 131618 79960
rect 130818 78752 131618 78872
rect 130818 77800 131618 77920
rect 130818 76848 131618 76968
rect 130818 75760 131618 75880
rect 130818 74808 131618 74928
rect 130818 73856 131618 73976
rect 130818 72768 131618 72888
rect 130818 71816 131618 71936
rect 130818 70864 131618 70984
rect 130818 69912 131618 70032
rect 130818 68824 131618 68944
rect 130818 67872 131618 67992
rect 130818 66920 131618 67040
rect 130818 65832 131618 65952
rect 130818 64880 131618 65000
rect 130818 63928 131618 64048
rect 130818 62840 131618 62960
rect 130818 61888 131618 62008
rect 130818 60936 131618 61056
rect 130818 59984 131618 60104
rect 130818 58896 131618 59016
rect 130818 57944 131618 58064
rect 130818 56992 131618 57112
rect 130818 55904 131618 56024
rect 130818 54952 131618 55072
rect 130818 54000 131618 54120
rect 130818 52912 131618 53032
rect 130818 51960 131618 52080
rect 130818 51008 131618 51128
rect 130818 50056 131618 50176
rect 130818 48968 131618 49088
rect 130818 48016 131618 48136
rect 130818 47064 131618 47184
rect 130818 45976 131618 46096
rect 130818 45024 131618 45144
rect 130818 44072 131618 44192
rect 130818 42984 131618 43104
rect 130818 42032 131618 42152
rect 130818 41080 131618 41200
rect 130818 40128 131618 40248
rect 130818 39040 131618 39160
rect 130818 38088 131618 38208
rect 130818 37136 131618 37256
rect 130818 36048 131618 36168
rect 130818 35096 131618 35216
rect 130818 34144 131618 34264
rect 130818 33056 131618 33176
rect 130818 32104 131618 32224
rect 130818 31152 131618 31272
rect 130818 30200 131618 30320
rect 130818 29112 131618 29232
rect 130818 28160 131618 28280
rect 130818 27208 131618 27328
rect 130818 26120 131618 26240
rect 130818 25168 131618 25288
rect 130818 24216 131618 24336
rect 130818 23128 131618 23248
rect 130818 22176 131618 22296
rect 130818 21224 131618 21344
rect 130818 20272 131618 20392
rect 130818 19184 131618 19304
rect 130818 18232 131618 18352
rect 130818 17280 131618 17400
rect 130818 16192 131618 16312
rect 130818 15240 131618 15360
rect 130818 14288 131618 14408
rect 130818 13200 131618 13320
rect 130818 12248 131618 12368
rect 130818 11296 131618 11416
rect 130818 10344 131618 10464
rect 130818 9256 131618 9376
rect 130818 8304 131618 8424
rect 130818 7352 131618 7472
rect 130818 6264 131618 6384
rect 130818 5312 131618 5432
rect 130818 4360 131618 4480
rect 130818 3272 131618 3392
rect 130818 2320 131618 2440
rect 130818 1368 131618 1488
rect 130818 416 131618 536
<< obsm3 >>
rect 735 129400 130738 129505
rect 735 128592 130818 129400
rect 735 128312 130738 128592
rect 735 127640 130818 128312
rect 735 127360 130738 127640
rect 735 126688 130818 127360
rect 735 126408 130738 126688
rect 735 125600 130818 126408
rect 735 125320 130738 125600
rect 735 124648 130818 125320
rect 735 124368 130738 124648
rect 735 123696 130818 124368
rect 735 123416 130738 123696
rect 735 122608 130818 123416
rect 735 122328 130738 122608
rect 735 121656 130818 122328
rect 735 121376 130738 121656
rect 735 120704 130818 121376
rect 735 120424 130738 120704
rect 735 119752 130818 120424
rect 735 119472 130738 119752
rect 735 118664 130818 119472
rect 735 118384 130738 118664
rect 735 117712 130818 118384
rect 735 117432 130738 117712
rect 735 116760 130818 117432
rect 735 116480 130738 116760
rect 735 115672 130818 116480
rect 735 115392 130738 115672
rect 735 114720 130818 115392
rect 735 114440 130738 114720
rect 735 113768 130818 114440
rect 735 113488 130738 113768
rect 735 112680 130818 113488
rect 735 112400 130738 112680
rect 735 111728 130818 112400
rect 735 111448 130738 111728
rect 735 110776 130818 111448
rect 735 110496 130738 110776
rect 735 109824 130818 110496
rect 735 109544 130738 109824
rect 735 108736 130818 109544
rect 735 108456 130738 108736
rect 735 107784 130818 108456
rect 735 107504 130738 107784
rect 735 106832 130818 107504
rect 735 106552 130738 106832
rect 735 105744 130818 106552
rect 735 105464 130738 105744
rect 735 104792 130818 105464
rect 735 104512 130738 104792
rect 735 103840 130818 104512
rect 735 103560 130738 103840
rect 735 102752 130818 103560
rect 735 102472 130738 102752
rect 735 101800 130818 102472
rect 735 101520 130738 101800
rect 735 100848 130818 101520
rect 735 100568 130738 100848
rect 735 99896 130818 100568
rect 735 99616 130738 99896
rect 735 98808 130818 99616
rect 735 98528 130738 98808
rect 735 97856 130818 98528
rect 735 97576 130738 97856
rect 735 96904 130818 97576
rect 735 96624 130738 96904
rect 735 95816 130818 96624
rect 735 95536 130738 95816
rect 735 94864 130818 95536
rect 735 94584 130738 94864
rect 735 93912 130818 94584
rect 735 93632 130738 93912
rect 735 92824 130818 93632
rect 735 92544 130738 92824
rect 735 91872 130818 92544
rect 735 91592 130738 91872
rect 735 90920 130818 91592
rect 735 90640 130738 90920
rect 735 89968 130818 90640
rect 735 89688 130738 89968
rect 735 88880 130818 89688
rect 735 88600 130738 88880
rect 735 87928 130818 88600
rect 735 87648 130738 87928
rect 735 86976 130818 87648
rect 735 86696 130738 86976
rect 735 85888 130818 86696
rect 735 85608 130738 85888
rect 735 84936 130818 85608
rect 735 84656 130738 84936
rect 735 83984 130818 84656
rect 735 83704 130738 83984
rect 735 82896 130818 83704
rect 735 82616 130738 82896
rect 735 81944 130818 82616
rect 735 81664 130738 81944
rect 735 80992 130818 81664
rect 735 80712 130738 80992
rect 735 80040 130818 80712
rect 735 79760 130738 80040
rect 735 78952 130818 79760
rect 735 78672 130738 78952
rect 735 78000 130818 78672
rect 735 77720 130738 78000
rect 735 77048 130818 77720
rect 735 76768 130738 77048
rect 735 75960 130818 76768
rect 735 75680 130738 75960
rect 735 75008 130818 75680
rect 735 74728 130738 75008
rect 735 74056 130818 74728
rect 735 73776 130738 74056
rect 735 72968 130818 73776
rect 735 72688 130738 72968
rect 735 72016 130818 72688
rect 735 71736 130738 72016
rect 735 71064 130818 71736
rect 735 70784 130738 71064
rect 735 70112 130818 70784
rect 735 69832 130738 70112
rect 735 69024 130818 69832
rect 735 68744 130738 69024
rect 735 68072 130818 68744
rect 735 67792 130738 68072
rect 735 67120 130818 67792
rect 735 66840 130738 67120
rect 735 66032 130818 66840
rect 735 65752 130738 66032
rect 735 65080 130818 65752
rect 735 64800 130738 65080
rect 735 64128 130818 64800
rect 735 63848 130738 64128
rect 735 63040 130818 63848
rect 735 62760 130738 63040
rect 735 62088 130818 62760
rect 735 61808 130738 62088
rect 735 61136 130818 61808
rect 735 60856 130738 61136
rect 735 60184 130818 60856
rect 735 59904 130738 60184
rect 735 59096 130818 59904
rect 735 58816 130738 59096
rect 735 58144 130818 58816
rect 735 57864 130738 58144
rect 735 57192 130818 57864
rect 735 56912 130738 57192
rect 735 56104 130818 56912
rect 735 55824 130738 56104
rect 735 55152 130818 55824
rect 735 54872 130738 55152
rect 735 54200 130818 54872
rect 735 53920 130738 54200
rect 735 53112 130818 53920
rect 735 52832 130738 53112
rect 735 52160 130818 52832
rect 735 51880 130738 52160
rect 735 51208 130818 51880
rect 735 50928 130738 51208
rect 735 50256 130818 50928
rect 735 49976 130738 50256
rect 735 49168 130818 49976
rect 735 48888 130738 49168
rect 735 48216 130818 48888
rect 735 47936 130738 48216
rect 735 47264 130818 47936
rect 735 46984 130738 47264
rect 735 46176 130818 46984
rect 735 45896 130738 46176
rect 735 45224 130818 45896
rect 735 44944 130738 45224
rect 735 44272 130818 44944
rect 735 43992 130738 44272
rect 735 43184 130818 43992
rect 735 42904 130738 43184
rect 735 42232 130818 42904
rect 735 41952 130738 42232
rect 735 41280 130818 41952
rect 735 41000 130738 41280
rect 735 40328 130818 41000
rect 735 40048 130738 40328
rect 735 39240 130818 40048
rect 735 38960 130738 39240
rect 735 38288 130818 38960
rect 735 38008 130738 38288
rect 735 37336 130818 38008
rect 735 37056 130738 37336
rect 735 36248 130818 37056
rect 735 35968 130738 36248
rect 735 35296 130818 35968
rect 735 35016 130738 35296
rect 735 34344 130818 35016
rect 735 34064 130738 34344
rect 735 33256 130818 34064
rect 735 32976 130738 33256
rect 735 32304 130818 32976
rect 735 32024 130738 32304
rect 735 31352 130818 32024
rect 735 31072 130738 31352
rect 735 30400 130818 31072
rect 735 30120 130738 30400
rect 735 29312 130818 30120
rect 735 29032 130738 29312
rect 735 28360 130818 29032
rect 735 28080 130738 28360
rect 735 27408 130818 28080
rect 735 27128 130738 27408
rect 735 26320 130818 27128
rect 735 26040 130738 26320
rect 735 25368 130818 26040
rect 735 25088 130738 25368
rect 735 24416 130818 25088
rect 735 24136 130738 24416
rect 735 23328 130818 24136
rect 735 23048 130738 23328
rect 735 22376 130818 23048
rect 735 22096 130738 22376
rect 735 21424 130818 22096
rect 735 21144 130738 21424
rect 735 20472 130818 21144
rect 735 20192 130738 20472
rect 735 19384 130818 20192
rect 735 19104 130738 19384
rect 735 18432 130818 19104
rect 735 18152 130738 18432
rect 735 17480 130818 18152
rect 735 17200 130738 17480
rect 735 16392 130818 17200
rect 735 16112 130738 16392
rect 735 15440 130818 16112
rect 735 15160 130738 15440
rect 735 14488 130818 15160
rect 735 14208 130738 14488
rect 735 13400 130818 14208
rect 735 13120 130738 13400
rect 735 12448 130818 13120
rect 735 12168 130738 12448
rect 735 11496 130818 12168
rect 735 11216 130738 11496
rect 735 10544 130818 11216
rect 735 10264 130738 10544
rect 735 9456 130818 10264
rect 735 9176 130738 9456
rect 735 8504 130818 9176
rect 735 8224 130738 8504
rect 735 7552 130818 8224
rect 735 7272 130738 7552
rect 735 6464 130818 7272
rect 735 6184 130738 6464
rect 735 5512 130818 6184
rect 735 5232 130738 5512
rect 735 4560 130818 5232
rect 735 4280 130738 4560
rect 735 3472 130818 4280
rect 735 3192 130738 3472
rect 735 2520 130818 3192
rect 735 2240 130738 2520
rect 735 1568 130818 2240
rect 735 1288 130738 1568
rect 735 616 130818 1288
rect 735 443 130738 616
<< metal4 >>
rect 3826 2128 4146 129520
rect 4486 2176 4806 129472
rect 5146 2176 5466 129472
rect 5806 2176 6126 129472
rect 19186 2128 19506 129520
rect 19846 2176 20166 129472
rect 20506 2176 20826 129472
rect 21166 2176 21486 129472
rect 34546 2128 34866 129520
rect 35206 2176 35526 129472
rect 35866 2176 36186 129472
rect 36526 2176 36846 129472
rect 49906 2128 50226 129520
rect 50566 2176 50886 129472
rect 51226 2176 51546 129472
rect 51886 2176 52206 129472
rect 65266 2128 65586 129520
rect 65926 2176 66246 129472
rect 66586 2176 66906 129472
rect 67246 2176 67566 129472
rect 80626 2128 80946 129520
rect 81286 2176 81606 129472
rect 81946 2176 82266 129472
rect 82606 2176 82926 129472
rect 95986 2128 96306 129520
rect 96646 2176 96966 129472
rect 97306 2176 97626 129472
rect 97966 2176 98286 129472
rect 111346 2128 111666 129520
rect 112006 2176 112326 129472
rect 112666 2176 112986 129472
rect 113326 2176 113646 129472
rect 126706 2128 127026 129520
rect 127366 2176 127686 129472
rect 128026 2176 128346 129472
rect 128686 2176 129006 129472
<< obsm4 >>
rect 9061 2619 19106 128485
rect 19586 2619 19766 128485
rect 20246 2619 20426 128485
rect 20906 2619 21086 128485
rect 21566 2619 34466 128485
rect 34946 2619 35126 128485
rect 35606 2619 35786 128485
rect 36266 2619 36446 128485
rect 36926 2619 49826 128485
rect 50306 2619 50486 128485
rect 50966 2619 51146 128485
rect 51626 2619 51806 128485
rect 52286 2619 65186 128485
rect 65666 2619 65846 128485
rect 66326 2619 66506 128485
rect 66986 2619 67166 128485
rect 67646 2619 80546 128485
rect 81026 2619 81206 128485
rect 81686 2619 81866 128485
rect 82346 2619 82526 128485
rect 83006 2619 95906 128485
rect 96386 2619 96566 128485
rect 97046 2619 97226 128485
rect 97706 2619 97886 128485
rect 98366 2619 111266 128485
rect 111746 2619 111926 128485
rect 112406 2619 112586 128485
rect 113066 2619 113246 128485
rect 113726 2619 126626 128485
rect 127106 2619 127255 128485
<< labels >>
rlabel metal3 s 130818 416 131618 536 6 clk
port 1 nsew signal input
rlabel metal2 s 128896 0 128952 800 6 flush_in
port 2 nsew signal input
rlabel metal2 s 4 0 60 800 6 i_in[0]
port 3 nsew signal input
rlabel metal2 s 7548 0 7604 800 6 i_in[10]
port 4 nsew signal input
rlabel metal2 s 8376 0 8432 800 6 i_in[11]
port 5 nsew signal input
rlabel metal2 s 9112 0 9168 800 6 i_in[12]
port 6 nsew signal input
rlabel metal2 s 9848 0 9904 800 6 i_in[13]
port 7 nsew signal input
rlabel metal2 s 10676 0 10732 800 6 i_in[14]
port 8 nsew signal input
rlabel metal2 s 11412 0 11468 800 6 i_in[15]
port 9 nsew signal input
rlabel metal2 s 12148 0 12204 800 6 i_in[16]
port 10 nsew signal input
rlabel metal2 s 12976 0 13032 800 6 i_in[17]
port 11 nsew signal input
rlabel metal2 s 13712 0 13768 800 6 i_in[18]
port 12 nsew signal input
rlabel metal2 s 14448 0 14504 800 6 i_in[19]
port 13 nsew signal input
rlabel metal2 s 740 0 796 800 6 i_in[1]
port 14 nsew signal input
rlabel metal2 s 15184 0 15240 800 6 i_in[20]
port 15 nsew signal input
rlabel metal2 s 16012 0 16068 800 6 i_in[21]
port 16 nsew signal input
rlabel metal2 s 16748 0 16804 800 6 i_in[22]
port 17 nsew signal input
rlabel metal2 s 17484 0 17540 800 6 i_in[23]
port 18 nsew signal input
rlabel metal2 s 18312 0 18368 800 6 i_in[24]
port 19 nsew signal input
rlabel metal2 s 19048 0 19104 800 6 i_in[25]
port 20 nsew signal input
rlabel metal2 s 19784 0 19840 800 6 i_in[26]
port 21 nsew signal input
rlabel metal2 s 20520 0 20576 800 6 i_in[27]
port 22 nsew signal input
rlabel metal2 s 21348 0 21404 800 6 i_in[28]
port 23 nsew signal input
rlabel metal2 s 22084 0 22140 800 6 i_in[29]
port 24 nsew signal input
rlabel metal2 s 1476 0 1532 800 6 i_in[2]
port 25 nsew signal input
rlabel metal2 s 22820 0 22876 800 6 i_in[30]
port 26 nsew signal input
rlabel metal2 s 23648 0 23704 800 6 i_in[31]
port 27 nsew signal input
rlabel metal2 s 24384 0 24440 800 6 i_in[32]
port 28 nsew signal input
rlabel metal2 s 25120 0 25176 800 6 i_in[33]
port 29 nsew signal input
rlabel metal2 s 25948 0 26004 800 6 i_in[34]
port 30 nsew signal input
rlabel metal2 s 26684 0 26740 800 6 i_in[35]
port 31 nsew signal input
rlabel metal2 s 27420 0 27476 800 6 i_in[36]
port 32 nsew signal input
rlabel metal2 s 28156 0 28212 800 6 i_in[37]
port 33 nsew signal input
rlabel metal2 s 28984 0 29040 800 6 i_in[38]
port 34 nsew signal input
rlabel metal2 s 29720 0 29776 800 6 i_in[39]
port 35 nsew signal input
rlabel metal2 s 2212 0 2268 800 6 i_in[3]
port 36 nsew signal input
rlabel metal2 s 30456 0 30512 800 6 i_in[40]
port 37 nsew signal input
rlabel metal2 s 31284 0 31340 800 6 i_in[41]
port 38 nsew signal input
rlabel metal2 s 32020 0 32076 800 6 i_in[42]
port 39 nsew signal input
rlabel metal2 s 32756 0 32812 800 6 i_in[43]
port 40 nsew signal input
rlabel metal2 s 33492 0 33548 800 6 i_in[44]
port 41 nsew signal input
rlabel metal2 s 34320 0 34376 800 6 i_in[45]
port 42 nsew signal input
rlabel metal2 s 35056 0 35112 800 6 i_in[46]
port 43 nsew signal input
rlabel metal2 s 35792 0 35848 800 6 i_in[47]
port 44 nsew signal input
rlabel metal2 s 36620 0 36676 800 6 i_in[48]
port 45 nsew signal input
rlabel metal2 s 37356 0 37412 800 6 i_in[49]
port 46 nsew signal input
rlabel metal2 s 3040 0 3096 800 6 i_in[4]
port 47 nsew signal input
rlabel metal2 s 38092 0 38148 800 6 i_in[50]
port 48 nsew signal input
rlabel metal2 s 38920 0 38976 800 6 i_in[51]
port 49 nsew signal input
rlabel metal2 s 39656 0 39712 800 6 i_in[52]
port 50 nsew signal input
rlabel metal2 s 40392 0 40448 800 6 i_in[53]
port 51 nsew signal input
rlabel metal2 s 41128 0 41184 800 6 i_in[54]
port 52 nsew signal input
rlabel metal2 s 41956 0 42012 800 6 i_in[55]
port 53 nsew signal input
rlabel metal2 s 42692 0 42748 800 6 i_in[56]
port 54 nsew signal input
rlabel metal2 s 43428 0 43484 800 6 i_in[57]
port 55 nsew signal input
rlabel metal2 s 44256 0 44312 800 6 i_in[58]
port 56 nsew signal input
rlabel metal2 s 44992 0 45048 800 6 i_in[59]
port 57 nsew signal input
rlabel metal2 s 3776 0 3832 800 6 i_in[5]
port 58 nsew signal input
rlabel metal2 s 45728 0 45784 800 6 i_in[60]
port 59 nsew signal input
rlabel metal2 s 46464 0 46520 800 6 i_in[61]
port 60 nsew signal input
rlabel metal2 s 47292 0 47348 800 6 i_in[62]
port 61 nsew signal input
rlabel metal2 s 48028 0 48084 800 6 i_in[63]
port 62 nsew signal input
rlabel metal2 s 48764 0 48820 800 6 i_in[64]
port 63 nsew signal input
rlabel metal2 s 49592 0 49648 800 6 i_in[65]
port 64 nsew signal input
rlabel metal2 s 50328 0 50384 800 6 i_in[66]
port 65 nsew signal input
rlabel metal2 s 51064 0 51120 800 6 i_in[67]
port 66 nsew signal input
rlabel metal2 s 51892 0 51948 800 6 i_in[68]
port 67 nsew signal input
rlabel metal2 s 52628 0 52684 800 6 i_in[69]
port 68 nsew signal input
rlabel metal2 s 4512 0 4568 800 6 i_in[6]
port 69 nsew signal input
rlabel metal2 s 5340 0 5396 800 6 i_in[7]
port 70 nsew signal input
rlabel metal2 s 6076 0 6132 800 6 i_in[8]
port 71 nsew signal input
rlabel metal2 s 6812 0 6868 800 6 i_in[9]
port 72 nsew signal input
rlabel metal2 s 53364 0 53420 800 6 i_out[0]
port 73 nsew signal output
rlabel metal2 s 61000 0 61056 800 6 i_out[10]
port 74 nsew signal output
rlabel metal2 s 61736 0 61792 800 6 i_out[11]
port 75 nsew signal output
rlabel metal2 s 62564 0 62620 800 6 i_out[12]
port 76 nsew signal output
rlabel metal2 s 63300 0 63356 800 6 i_out[13]
port 77 nsew signal output
rlabel metal2 s 64036 0 64092 800 6 i_out[14]
port 78 nsew signal output
rlabel metal2 s 64864 0 64920 800 6 i_out[15]
port 79 nsew signal output
rlabel metal2 s 65600 0 65656 800 6 i_out[16]
port 80 nsew signal output
rlabel metal2 s 66336 0 66392 800 6 i_out[17]
port 81 nsew signal output
rlabel metal2 s 67072 0 67128 800 6 i_out[18]
port 82 nsew signal output
rlabel metal2 s 67900 0 67956 800 6 i_out[19]
port 83 nsew signal output
rlabel metal2 s 54100 0 54156 800 6 i_out[1]
port 84 nsew signal output
rlabel metal2 s 68636 0 68692 800 6 i_out[20]
port 85 nsew signal output
rlabel metal2 s 69372 0 69428 800 6 i_out[21]
port 86 nsew signal output
rlabel metal2 s 70200 0 70256 800 6 i_out[22]
port 87 nsew signal output
rlabel metal2 s 70936 0 70992 800 6 i_out[23]
port 88 nsew signal output
rlabel metal2 s 71672 0 71728 800 6 i_out[24]
port 89 nsew signal output
rlabel metal2 s 72500 0 72556 800 6 i_out[25]
port 90 nsew signal output
rlabel metal2 s 73236 0 73292 800 6 i_out[26]
port 91 nsew signal output
rlabel metal2 s 73972 0 74028 800 6 i_out[27]
port 92 nsew signal output
rlabel metal2 s 74708 0 74764 800 6 i_out[28]
port 93 nsew signal output
rlabel metal2 s 75536 0 75592 800 6 i_out[29]
port 94 nsew signal output
rlabel metal2 s 54928 0 54984 800 6 i_out[2]
port 95 nsew signal output
rlabel metal2 s 76272 0 76328 800 6 i_out[30]
port 96 nsew signal output
rlabel metal2 s 77008 0 77064 800 6 i_out[31]
port 97 nsew signal output
rlabel metal2 s 77836 0 77892 800 6 i_out[32]
port 98 nsew signal output
rlabel metal2 s 78572 0 78628 800 6 i_out[33]
port 99 nsew signal output
rlabel metal2 s 79308 0 79364 800 6 i_out[34]
port 100 nsew signal output
rlabel metal2 s 80044 0 80100 800 6 i_out[35]
port 101 nsew signal output
rlabel metal2 s 80872 0 80928 800 6 i_out[36]
port 102 nsew signal output
rlabel metal2 s 81608 0 81664 800 6 i_out[37]
port 103 nsew signal output
rlabel metal2 s 82344 0 82400 800 6 i_out[38]
port 104 nsew signal output
rlabel metal2 s 83172 0 83228 800 6 i_out[39]
port 105 nsew signal output
rlabel metal2 s 55664 0 55720 800 6 i_out[3]
port 106 nsew signal output
rlabel metal2 s 83908 0 83964 800 6 i_out[40]
port 107 nsew signal output
rlabel metal2 s 84644 0 84700 800 6 i_out[41]
port 108 nsew signal output
rlabel metal2 s 85472 0 85528 800 6 i_out[42]
port 109 nsew signal output
rlabel metal2 s 86208 0 86264 800 6 i_out[43]
port 110 nsew signal output
rlabel metal2 s 86944 0 87000 800 6 i_out[44]
port 111 nsew signal output
rlabel metal2 s 87680 0 87736 800 6 i_out[45]
port 112 nsew signal output
rlabel metal2 s 88508 0 88564 800 6 i_out[46]
port 113 nsew signal output
rlabel metal2 s 89244 0 89300 800 6 i_out[47]
port 114 nsew signal output
rlabel metal2 s 89980 0 90036 800 6 i_out[48]
port 115 nsew signal output
rlabel metal2 s 90808 0 90864 800 6 i_out[49]
port 116 nsew signal output
rlabel metal2 s 56400 0 56456 800 6 i_out[4]
port 117 nsew signal output
rlabel metal2 s 91544 0 91600 800 6 i_out[50]
port 118 nsew signal output
rlabel metal2 s 92280 0 92336 800 6 i_out[51]
port 119 nsew signal output
rlabel metal2 s 93016 0 93072 800 6 i_out[52]
port 120 nsew signal output
rlabel metal2 s 93844 0 93900 800 6 i_out[53]
port 121 nsew signal output
rlabel metal2 s 94580 0 94636 800 6 i_out[54]
port 122 nsew signal output
rlabel metal2 s 95316 0 95372 800 6 i_out[55]
port 123 nsew signal output
rlabel metal2 s 96144 0 96200 800 6 i_out[56]
port 124 nsew signal output
rlabel metal2 s 96880 0 96936 800 6 i_out[57]
port 125 nsew signal output
rlabel metal2 s 97616 0 97672 800 6 i_out[58]
port 126 nsew signal output
rlabel metal2 s 98444 0 98500 800 6 i_out[59]
port 127 nsew signal output
rlabel metal2 s 57228 0 57284 800 6 i_out[5]
port 128 nsew signal output
rlabel metal2 s 99180 0 99236 800 6 i_out[60]
port 129 nsew signal output
rlabel metal2 s 99916 0 99972 800 6 i_out[61]
port 130 nsew signal output
rlabel metal2 s 100652 0 100708 800 6 i_out[62]
port 131 nsew signal output
rlabel metal2 s 101480 0 101536 800 6 i_out[63]
port 132 nsew signal output
rlabel metal2 s 102216 0 102272 800 6 i_out[64]
port 133 nsew signal output
rlabel metal2 s 102952 0 103008 800 6 i_out[65]
port 134 nsew signal output
rlabel metal2 s 103780 0 103836 800 6 i_out[66]
port 135 nsew signal output
rlabel metal2 s 104516 0 104572 800 6 i_out[67]
port 136 nsew signal output
rlabel metal2 s 105252 0 105308 800 6 i_out[68]
port 137 nsew signal output
rlabel metal2 s 105988 0 106044 800 6 i_out[69]
port 138 nsew signal output
rlabel metal2 s 57964 0 58020 800 6 i_out[6]
port 139 nsew signal output
rlabel metal2 s 106816 0 106872 800 6 i_out[70]
port 140 nsew signal output
rlabel metal2 s 107552 0 107608 800 6 i_out[71]
port 141 nsew signal output
rlabel metal2 s 108288 0 108344 800 6 i_out[72]
port 142 nsew signal output
rlabel metal2 s 109116 0 109172 800 6 i_out[73]
port 143 nsew signal output
rlabel metal2 s 109852 0 109908 800 6 i_out[74]
port 144 nsew signal output
rlabel metal2 s 110588 0 110644 800 6 i_out[75]
port 145 nsew signal output
rlabel metal2 s 111416 0 111472 800 6 i_out[76]
port 146 nsew signal output
rlabel metal2 s 112152 0 112208 800 6 i_out[77]
port 147 nsew signal output
rlabel metal2 s 112888 0 112944 800 6 i_out[78]
port 148 nsew signal output
rlabel metal2 s 113624 0 113680 800 6 i_out[79]
port 149 nsew signal output
rlabel metal2 s 58700 0 58756 800 6 i_out[7]
port 150 nsew signal output
rlabel metal2 s 114452 0 114508 800 6 i_out[80]
port 151 nsew signal output
rlabel metal2 s 115188 0 115244 800 6 i_out[81]
port 152 nsew signal output
rlabel metal2 s 115924 0 115980 800 6 i_out[82]
port 153 nsew signal output
rlabel metal2 s 116752 0 116808 800 6 i_out[83]
port 154 nsew signal output
rlabel metal2 s 117488 0 117544 800 6 i_out[84]
port 155 nsew signal output
rlabel metal2 s 118224 0 118280 800 6 i_out[85]
port 156 nsew signal output
rlabel metal2 s 118960 0 119016 800 6 i_out[86]
port 157 nsew signal output
rlabel metal2 s 119788 0 119844 800 6 i_out[87]
port 158 nsew signal output
rlabel metal2 s 120524 0 120580 800 6 i_out[88]
port 159 nsew signal output
rlabel metal2 s 121260 0 121316 800 6 i_out[89]
port 160 nsew signal output
rlabel metal2 s 59436 0 59492 800 6 i_out[8]
port 161 nsew signal output
rlabel metal2 s 122088 0 122144 800 6 i_out[90]
port 162 nsew signal output
rlabel metal2 s 122824 0 122880 800 6 i_out[91]
port 163 nsew signal output
rlabel metal2 s 123560 0 123616 800 6 i_out[92]
port 164 nsew signal output
rlabel metal2 s 124388 0 124444 800 6 i_out[93]
port 165 nsew signal output
rlabel metal2 s 125124 0 125180 800 6 i_out[94]
port 166 nsew signal output
rlabel metal2 s 125860 0 125916 800 6 i_out[95]
port 167 nsew signal output
rlabel metal2 s 126596 0 126652 800 6 i_out[96]
port 168 nsew signal output
rlabel metal2 s 127424 0 127480 800 6 i_out[97]
port 169 nsew signal output
rlabel metal2 s 128160 0 128216 800 6 i_out[98]
port 170 nsew signal output
rlabel metal2 s 60264 0 60320 800 6 i_out[9]
port 171 nsew signal output
rlabel metal2 s 129724 0 129780 800 6 inval_in
port 172 nsew signal input
rlabel metal3 s 130818 2320 131618 2440 6 m_in[0]
port 173 nsew signal input
rlabel metal3 s 130818 101600 131618 101720 6 m_in[100]
port 174 nsew signal input
rlabel metal3 s 130818 102552 131618 102672 6 m_in[101]
port 175 nsew signal input
rlabel metal3 s 130818 103640 131618 103760 6 m_in[102]
port 176 nsew signal input
rlabel metal3 s 130818 104592 131618 104712 6 m_in[103]
port 177 nsew signal input
rlabel metal3 s 130818 105544 131618 105664 6 m_in[104]
port 178 nsew signal input
rlabel metal3 s 130818 106632 131618 106752 6 m_in[105]
port 179 nsew signal input
rlabel metal3 s 130818 107584 131618 107704 6 m_in[106]
port 180 nsew signal input
rlabel metal3 s 130818 108536 131618 108656 6 m_in[107]
port 181 nsew signal input
rlabel metal3 s 130818 109624 131618 109744 6 m_in[108]
port 182 nsew signal input
rlabel metal3 s 130818 110576 131618 110696 6 m_in[109]
port 183 nsew signal input
rlabel metal3 s 130818 12248 131618 12368 6 m_in[10]
port 184 nsew signal input
rlabel metal3 s 130818 111528 131618 111648 6 m_in[110]
port 185 nsew signal input
rlabel metal3 s 130818 112480 131618 112600 6 m_in[111]
port 186 nsew signal input
rlabel metal3 s 130818 113568 131618 113688 6 m_in[112]
port 187 nsew signal input
rlabel metal3 s 130818 114520 131618 114640 6 m_in[113]
port 188 nsew signal input
rlabel metal3 s 130818 115472 131618 115592 6 m_in[114]
port 189 nsew signal input
rlabel metal3 s 130818 116560 131618 116680 6 m_in[115]
port 190 nsew signal input
rlabel metal3 s 130818 117512 131618 117632 6 m_in[116]
port 191 nsew signal input
rlabel metal3 s 130818 118464 131618 118584 6 m_in[117]
port 192 nsew signal input
rlabel metal3 s 130818 119552 131618 119672 6 m_in[118]
port 193 nsew signal input
rlabel metal3 s 130818 120504 131618 120624 6 m_in[119]
port 194 nsew signal input
rlabel metal3 s 130818 13200 131618 13320 6 m_in[11]
port 195 nsew signal input
rlabel metal3 s 130818 121456 131618 121576 6 m_in[120]
port 196 nsew signal input
rlabel metal3 s 130818 122408 131618 122528 6 m_in[121]
port 197 nsew signal input
rlabel metal3 s 130818 123496 131618 123616 6 m_in[122]
port 198 nsew signal input
rlabel metal3 s 130818 124448 131618 124568 6 m_in[123]
port 199 nsew signal input
rlabel metal3 s 130818 125400 131618 125520 6 m_in[124]
port 200 nsew signal input
rlabel metal3 s 130818 126488 131618 126608 6 m_in[125]
port 201 nsew signal input
rlabel metal3 s 130818 127440 131618 127560 6 m_in[126]
port 202 nsew signal input
rlabel metal3 s 130818 128392 131618 128512 6 m_in[127]
port 203 nsew signal input
rlabel metal3 s 130818 129480 131618 129600 6 m_in[128]
port 204 nsew signal input
rlabel metal3 s 130818 130432 131618 130552 6 m_in[129]
port 205 nsew signal input
rlabel metal3 s 130818 14288 131618 14408 6 m_in[12]
port 206 nsew signal input
rlabel metal3 s 130818 131384 131618 131504 6 m_in[130]
port 207 nsew signal input
rlabel metal3 s 130818 15240 131618 15360 6 m_in[13]
port 208 nsew signal input
rlabel metal3 s 130818 16192 131618 16312 6 m_in[14]
port 209 nsew signal input
rlabel metal3 s 130818 17280 131618 17400 6 m_in[15]
port 210 nsew signal input
rlabel metal3 s 130818 18232 131618 18352 6 m_in[16]
port 211 nsew signal input
rlabel metal3 s 130818 19184 131618 19304 6 m_in[17]
port 212 nsew signal input
rlabel metal3 s 130818 20272 131618 20392 6 m_in[18]
port 213 nsew signal input
rlabel metal3 s 130818 21224 131618 21344 6 m_in[19]
port 214 nsew signal input
rlabel metal3 s 130818 3272 131618 3392 6 m_in[1]
port 215 nsew signal input
rlabel metal3 s 130818 22176 131618 22296 6 m_in[20]
port 216 nsew signal input
rlabel metal3 s 130818 23128 131618 23248 6 m_in[21]
port 217 nsew signal input
rlabel metal3 s 130818 24216 131618 24336 6 m_in[22]
port 218 nsew signal input
rlabel metal3 s 130818 25168 131618 25288 6 m_in[23]
port 219 nsew signal input
rlabel metal3 s 130818 26120 131618 26240 6 m_in[24]
port 220 nsew signal input
rlabel metal3 s 130818 27208 131618 27328 6 m_in[25]
port 221 nsew signal input
rlabel metal3 s 130818 28160 131618 28280 6 m_in[26]
port 222 nsew signal input
rlabel metal3 s 130818 29112 131618 29232 6 m_in[27]
port 223 nsew signal input
rlabel metal3 s 130818 30200 131618 30320 6 m_in[28]
port 224 nsew signal input
rlabel metal3 s 130818 31152 131618 31272 6 m_in[29]
port 225 nsew signal input
rlabel metal3 s 130818 4360 131618 4480 6 m_in[2]
port 226 nsew signal input
rlabel metal3 s 130818 32104 131618 32224 6 m_in[30]
port 227 nsew signal input
rlabel metal3 s 130818 33056 131618 33176 6 m_in[31]
port 228 nsew signal input
rlabel metal3 s 130818 34144 131618 34264 6 m_in[32]
port 229 nsew signal input
rlabel metal3 s 130818 35096 131618 35216 6 m_in[33]
port 230 nsew signal input
rlabel metal3 s 130818 36048 131618 36168 6 m_in[34]
port 231 nsew signal input
rlabel metal3 s 130818 37136 131618 37256 6 m_in[35]
port 232 nsew signal input
rlabel metal3 s 130818 38088 131618 38208 6 m_in[36]
port 233 nsew signal input
rlabel metal3 s 130818 39040 131618 39160 6 m_in[37]
port 234 nsew signal input
rlabel metal3 s 130818 40128 131618 40248 6 m_in[38]
port 235 nsew signal input
rlabel metal3 s 130818 41080 131618 41200 6 m_in[39]
port 236 nsew signal input
rlabel metal3 s 130818 5312 131618 5432 6 m_in[3]
port 237 nsew signal input
rlabel metal3 s 130818 42032 131618 42152 6 m_in[40]
port 238 nsew signal input
rlabel metal3 s 130818 42984 131618 43104 6 m_in[41]
port 239 nsew signal input
rlabel metal3 s 130818 44072 131618 44192 6 m_in[42]
port 240 nsew signal input
rlabel metal3 s 130818 45024 131618 45144 6 m_in[43]
port 241 nsew signal input
rlabel metal3 s 130818 45976 131618 46096 6 m_in[44]
port 242 nsew signal input
rlabel metal3 s 130818 47064 131618 47184 6 m_in[45]
port 243 nsew signal input
rlabel metal3 s 130818 48016 131618 48136 6 m_in[46]
port 244 nsew signal input
rlabel metal3 s 130818 48968 131618 49088 6 m_in[47]
port 245 nsew signal input
rlabel metal3 s 130818 50056 131618 50176 6 m_in[48]
port 246 nsew signal input
rlabel metal3 s 130818 51008 131618 51128 6 m_in[49]
port 247 nsew signal input
rlabel metal3 s 130818 6264 131618 6384 6 m_in[4]
port 248 nsew signal input
rlabel metal3 s 130818 51960 131618 52080 6 m_in[50]
port 249 nsew signal input
rlabel metal3 s 130818 52912 131618 53032 6 m_in[51]
port 250 nsew signal input
rlabel metal3 s 130818 54000 131618 54120 6 m_in[52]
port 251 nsew signal input
rlabel metal3 s 130818 54952 131618 55072 6 m_in[53]
port 252 nsew signal input
rlabel metal3 s 130818 55904 131618 56024 6 m_in[54]
port 253 nsew signal input
rlabel metal3 s 130818 56992 131618 57112 6 m_in[55]
port 254 nsew signal input
rlabel metal3 s 130818 57944 131618 58064 6 m_in[56]
port 255 nsew signal input
rlabel metal3 s 130818 58896 131618 59016 6 m_in[57]
port 256 nsew signal input
rlabel metal3 s 130818 59984 131618 60104 6 m_in[58]
port 257 nsew signal input
rlabel metal3 s 130818 60936 131618 61056 6 m_in[59]
port 258 nsew signal input
rlabel metal3 s 130818 7352 131618 7472 6 m_in[5]
port 259 nsew signal input
rlabel metal3 s 130818 61888 131618 62008 6 m_in[60]
port 260 nsew signal input
rlabel metal3 s 130818 62840 131618 62960 6 m_in[61]
port 261 nsew signal input
rlabel metal3 s 130818 63928 131618 64048 6 m_in[62]
port 262 nsew signal input
rlabel metal3 s 130818 64880 131618 65000 6 m_in[63]
port 263 nsew signal input
rlabel metal3 s 130818 65832 131618 65952 6 m_in[64]
port 264 nsew signal input
rlabel metal3 s 130818 66920 131618 67040 6 m_in[65]
port 265 nsew signal input
rlabel metal3 s 130818 67872 131618 67992 6 m_in[66]
port 266 nsew signal input
rlabel metal3 s 130818 68824 131618 68944 6 m_in[67]
port 267 nsew signal input
rlabel metal3 s 130818 69912 131618 70032 6 m_in[68]
port 268 nsew signal input
rlabel metal3 s 130818 70864 131618 70984 6 m_in[69]
port 269 nsew signal input
rlabel metal3 s 130818 8304 131618 8424 6 m_in[6]
port 270 nsew signal input
rlabel metal3 s 130818 71816 131618 71936 6 m_in[70]
port 271 nsew signal input
rlabel metal3 s 130818 72768 131618 72888 6 m_in[71]
port 272 nsew signal input
rlabel metal3 s 130818 73856 131618 73976 6 m_in[72]
port 273 nsew signal input
rlabel metal3 s 130818 74808 131618 74928 6 m_in[73]
port 274 nsew signal input
rlabel metal3 s 130818 75760 131618 75880 6 m_in[74]
port 275 nsew signal input
rlabel metal3 s 130818 76848 131618 76968 6 m_in[75]
port 276 nsew signal input
rlabel metal3 s 130818 77800 131618 77920 6 m_in[76]
port 277 nsew signal input
rlabel metal3 s 130818 78752 131618 78872 6 m_in[77]
port 278 nsew signal input
rlabel metal3 s 130818 79840 131618 79960 6 m_in[78]
port 279 nsew signal input
rlabel metal3 s 130818 80792 131618 80912 6 m_in[79]
port 280 nsew signal input
rlabel metal3 s 130818 9256 131618 9376 6 m_in[7]
port 281 nsew signal input
rlabel metal3 s 130818 81744 131618 81864 6 m_in[80]
port 282 nsew signal input
rlabel metal3 s 130818 82696 131618 82816 6 m_in[81]
port 283 nsew signal input
rlabel metal3 s 130818 83784 131618 83904 6 m_in[82]
port 284 nsew signal input
rlabel metal3 s 130818 84736 131618 84856 6 m_in[83]
port 285 nsew signal input
rlabel metal3 s 130818 85688 131618 85808 6 m_in[84]
port 286 nsew signal input
rlabel metal3 s 130818 86776 131618 86896 6 m_in[85]
port 287 nsew signal input
rlabel metal3 s 130818 87728 131618 87848 6 m_in[86]
port 288 nsew signal input
rlabel metal3 s 130818 88680 131618 88800 6 m_in[87]
port 289 nsew signal input
rlabel metal3 s 130818 89768 131618 89888 6 m_in[88]
port 290 nsew signal input
rlabel metal3 s 130818 90720 131618 90840 6 m_in[89]
port 291 nsew signal input
rlabel metal3 s 130818 10344 131618 10464 6 m_in[8]
port 292 nsew signal input
rlabel metal3 s 130818 91672 131618 91792 6 m_in[90]
port 293 nsew signal input
rlabel metal3 s 130818 92624 131618 92744 6 m_in[91]
port 294 nsew signal input
rlabel metal3 s 130818 93712 131618 93832 6 m_in[92]
port 295 nsew signal input
rlabel metal3 s 130818 94664 131618 94784 6 m_in[93]
port 296 nsew signal input
rlabel metal3 s 130818 95616 131618 95736 6 m_in[94]
port 297 nsew signal input
rlabel metal3 s 130818 96704 131618 96824 6 m_in[95]
port 298 nsew signal input
rlabel metal3 s 130818 97656 131618 97776 6 m_in[96]
port 299 nsew signal input
rlabel metal3 s 130818 98608 131618 98728 6 m_in[97]
port 300 nsew signal input
rlabel metal3 s 130818 99696 131618 99816 6 m_in[98]
port 301 nsew signal input
rlabel metal3 s 130818 100648 131618 100768 6 m_in[99]
port 302 nsew signal input
rlabel metal3 s 130818 11296 131618 11416 6 m_in[9]
port 303 nsew signal input
rlabel metal3 s 130818 1368 131618 1488 6 rst
port 304 nsew signal input
rlabel metal2 s 130460 0 130516 800 6 stall_in
port 305 nsew signal input
rlabel metal2 s 131196 0 131252 800 6 stall_out
port 306 nsew signal output
rlabel metal2 s 4 131200 60 132000 6 wishbone_in[0]
port 307 nsew signal input
rlabel metal2 s 7548 131200 7604 132000 6 wishbone_in[10]
port 308 nsew signal input
rlabel metal2 s 8376 131200 8432 132000 6 wishbone_in[11]
port 309 nsew signal input
rlabel metal2 s 9112 131200 9168 132000 6 wishbone_in[12]
port 310 nsew signal input
rlabel metal2 s 9848 131200 9904 132000 6 wishbone_in[13]
port 311 nsew signal input
rlabel metal2 s 10676 131200 10732 132000 6 wishbone_in[14]
port 312 nsew signal input
rlabel metal2 s 11412 131200 11468 132000 6 wishbone_in[15]
port 313 nsew signal input
rlabel metal2 s 12148 131200 12204 132000 6 wishbone_in[16]
port 314 nsew signal input
rlabel metal2 s 12976 131200 13032 132000 6 wishbone_in[17]
port 315 nsew signal input
rlabel metal2 s 13712 131200 13768 132000 6 wishbone_in[18]
port 316 nsew signal input
rlabel metal2 s 14448 131200 14504 132000 6 wishbone_in[19]
port 317 nsew signal input
rlabel metal2 s 740 131200 796 132000 6 wishbone_in[1]
port 318 nsew signal input
rlabel metal2 s 15184 131200 15240 132000 6 wishbone_in[20]
port 319 nsew signal input
rlabel metal2 s 16012 131200 16068 132000 6 wishbone_in[21]
port 320 nsew signal input
rlabel metal2 s 16748 131200 16804 132000 6 wishbone_in[22]
port 321 nsew signal input
rlabel metal2 s 17484 131200 17540 132000 6 wishbone_in[23]
port 322 nsew signal input
rlabel metal2 s 18312 131200 18368 132000 6 wishbone_in[24]
port 323 nsew signal input
rlabel metal2 s 19048 131200 19104 132000 6 wishbone_in[25]
port 324 nsew signal input
rlabel metal2 s 19784 131200 19840 132000 6 wishbone_in[26]
port 325 nsew signal input
rlabel metal2 s 20520 131200 20576 132000 6 wishbone_in[27]
port 326 nsew signal input
rlabel metal2 s 21348 131200 21404 132000 6 wishbone_in[28]
port 327 nsew signal input
rlabel metal2 s 22084 131200 22140 132000 6 wishbone_in[29]
port 328 nsew signal input
rlabel metal2 s 1476 131200 1532 132000 6 wishbone_in[2]
port 329 nsew signal input
rlabel metal2 s 22820 131200 22876 132000 6 wishbone_in[30]
port 330 nsew signal input
rlabel metal2 s 23648 131200 23704 132000 6 wishbone_in[31]
port 331 nsew signal input
rlabel metal2 s 24384 131200 24440 132000 6 wishbone_in[32]
port 332 nsew signal input
rlabel metal2 s 25120 131200 25176 132000 6 wishbone_in[33]
port 333 nsew signal input
rlabel metal2 s 25948 131200 26004 132000 6 wishbone_in[34]
port 334 nsew signal input
rlabel metal2 s 26684 131200 26740 132000 6 wishbone_in[35]
port 335 nsew signal input
rlabel metal2 s 27420 131200 27476 132000 6 wishbone_in[36]
port 336 nsew signal input
rlabel metal2 s 28156 131200 28212 132000 6 wishbone_in[37]
port 337 nsew signal input
rlabel metal2 s 28984 131200 29040 132000 6 wishbone_in[38]
port 338 nsew signal input
rlabel metal2 s 29720 131200 29776 132000 6 wishbone_in[39]
port 339 nsew signal input
rlabel metal2 s 2212 131200 2268 132000 6 wishbone_in[3]
port 340 nsew signal input
rlabel metal2 s 30456 131200 30512 132000 6 wishbone_in[40]
port 341 nsew signal input
rlabel metal2 s 31284 131200 31340 132000 6 wishbone_in[41]
port 342 nsew signal input
rlabel metal2 s 32020 131200 32076 132000 6 wishbone_in[42]
port 343 nsew signal input
rlabel metal2 s 32756 131200 32812 132000 6 wishbone_in[43]
port 344 nsew signal input
rlabel metal2 s 33492 131200 33548 132000 6 wishbone_in[44]
port 345 nsew signal input
rlabel metal2 s 34320 131200 34376 132000 6 wishbone_in[45]
port 346 nsew signal input
rlabel metal2 s 35056 131200 35112 132000 6 wishbone_in[46]
port 347 nsew signal input
rlabel metal2 s 35792 131200 35848 132000 6 wishbone_in[47]
port 348 nsew signal input
rlabel metal2 s 36620 131200 36676 132000 6 wishbone_in[48]
port 349 nsew signal input
rlabel metal2 s 37356 131200 37412 132000 6 wishbone_in[49]
port 350 nsew signal input
rlabel metal2 s 3040 131200 3096 132000 6 wishbone_in[4]
port 351 nsew signal input
rlabel metal2 s 38092 131200 38148 132000 6 wishbone_in[50]
port 352 nsew signal input
rlabel metal2 s 38920 131200 38976 132000 6 wishbone_in[51]
port 353 nsew signal input
rlabel metal2 s 39656 131200 39712 132000 6 wishbone_in[52]
port 354 nsew signal input
rlabel metal2 s 40392 131200 40448 132000 6 wishbone_in[53]
port 355 nsew signal input
rlabel metal2 s 41128 131200 41184 132000 6 wishbone_in[54]
port 356 nsew signal input
rlabel metal2 s 41956 131200 42012 132000 6 wishbone_in[55]
port 357 nsew signal input
rlabel metal2 s 42692 131200 42748 132000 6 wishbone_in[56]
port 358 nsew signal input
rlabel metal2 s 43428 131200 43484 132000 6 wishbone_in[57]
port 359 nsew signal input
rlabel metal2 s 44256 131200 44312 132000 6 wishbone_in[58]
port 360 nsew signal input
rlabel metal2 s 44992 131200 45048 132000 6 wishbone_in[59]
port 361 nsew signal input
rlabel metal2 s 3776 131200 3832 132000 6 wishbone_in[5]
port 362 nsew signal input
rlabel metal2 s 45728 131200 45784 132000 6 wishbone_in[60]
port 363 nsew signal input
rlabel metal2 s 46464 131200 46520 132000 6 wishbone_in[61]
port 364 nsew signal input
rlabel metal2 s 47292 131200 47348 132000 6 wishbone_in[62]
port 365 nsew signal input
rlabel metal2 s 48028 131200 48084 132000 6 wishbone_in[63]
port 366 nsew signal input
rlabel metal2 s 48764 131200 48820 132000 6 wishbone_in[64]
port 367 nsew signal input
rlabel metal2 s 49592 131200 49648 132000 6 wishbone_in[65]
port 368 nsew signal input
rlabel metal2 s 4512 131200 4568 132000 6 wishbone_in[6]
port 369 nsew signal input
rlabel metal2 s 5340 131200 5396 132000 6 wishbone_in[7]
port 370 nsew signal input
rlabel metal2 s 6076 131200 6132 132000 6 wishbone_in[8]
port 371 nsew signal input
rlabel metal2 s 6812 131200 6868 132000 6 wishbone_in[9]
port 372 nsew signal input
rlabel metal2 s 50328 131200 50384 132000 6 wishbone_out[0]
port 373 nsew signal output
rlabel metal2 s 126596 131200 126652 132000 6 wishbone_out[100]
port 374 nsew signal output
rlabel metal2 s 127424 131200 127480 132000 6 wishbone_out[101]
port 375 nsew signal output
rlabel metal2 s 128160 131200 128216 132000 6 wishbone_out[102]
port 376 nsew signal output
rlabel metal2 s 128896 131200 128952 132000 6 wishbone_out[103]
port 377 nsew signal output
rlabel metal2 s 129724 131200 129780 132000 6 wishbone_out[104]
port 378 nsew signal output
rlabel metal2 s 130460 131200 130516 132000 6 wishbone_out[105]
port 379 nsew signal output
rlabel metal2 s 131196 131200 131252 132000 6 wishbone_out[106]
port 380 nsew signal output
rlabel metal2 s 57964 131200 58020 132000 6 wishbone_out[10]
port 381 nsew signal output
rlabel metal2 s 58700 131200 58756 132000 6 wishbone_out[11]
port 382 nsew signal output
rlabel metal2 s 59436 131200 59492 132000 6 wishbone_out[12]
port 383 nsew signal output
rlabel metal2 s 60264 131200 60320 132000 6 wishbone_out[13]
port 384 nsew signal output
rlabel metal2 s 61000 131200 61056 132000 6 wishbone_out[14]
port 385 nsew signal output
rlabel metal2 s 61736 131200 61792 132000 6 wishbone_out[15]
port 386 nsew signal output
rlabel metal2 s 62564 131200 62620 132000 6 wishbone_out[16]
port 387 nsew signal output
rlabel metal2 s 63300 131200 63356 132000 6 wishbone_out[17]
port 388 nsew signal output
rlabel metal2 s 64036 131200 64092 132000 6 wishbone_out[18]
port 389 nsew signal output
rlabel metal2 s 64864 131200 64920 132000 6 wishbone_out[19]
port 390 nsew signal output
rlabel metal2 s 51064 131200 51120 132000 6 wishbone_out[1]
port 391 nsew signal output
rlabel metal2 s 65600 131200 65656 132000 6 wishbone_out[20]
port 392 nsew signal output
rlabel metal2 s 66336 131200 66392 132000 6 wishbone_out[21]
port 393 nsew signal output
rlabel metal2 s 67072 131200 67128 132000 6 wishbone_out[22]
port 394 nsew signal output
rlabel metal2 s 67900 131200 67956 132000 6 wishbone_out[23]
port 395 nsew signal output
rlabel metal2 s 68636 131200 68692 132000 6 wishbone_out[24]
port 396 nsew signal output
rlabel metal2 s 69372 131200 69428 132000 6 wishbone_out[25]
port 397 nsew signal output
rlabel metal2 s 70200 131200 70256 132000 6 wishbone_out[26]
port 398 nsew signal output
rlabel metal2 s 70936 131200 70992 132000 6 wishbone_out[27]
port 399 nsew signal output
rlabel metal2 s 71672 131200 71728 132000 6 wishbone_out[28]
port 400 nsew signal output
rlabel metal2 s 72500 131200 72556 132000 6 wishbone_out[29]
port 401 nsew signal output
rlabel metal2 s 51892 131200 51948 132000 6 wishbone_out[2]
port 402 nsew signal output
rlabel metal2 s 73236 131200 73292 132000 6 wishbone_out[30]
port 403 nsew signal output
rlabel metal2 s 73972 131200 74028 132000 6 wishbone_out[31]
port 404 nsew signal output
rlabel metal2 s 74708 131200 74764 132000 6 wishbone_out[32]
port 405 nsew signal output
rlabel metal2 s 75536 131200 75592 132000 6 wishbone_out[33]
port 406 nsew signal output
rlabel metal2 s 76272 131200 76328 132000 6 wishbone_out[34]
port 407 nsew signal output
rlabel metal2 s 77008 131200 77064 132000 6 wishbone_out[35]
port 408 nsew signal output
rlabel metal2 s 77836 131200 77892 132000 6 wishbone_out[36]
port 409 nsew signal output
rlabel metal2 s 78572 131200 78628 132000 6 wishbone_out[37]
port 410 nsew signal output
rlabel metal2 s 79308 131200 79364 132000 6 wishbone_out[38]
port 411 nsew signal output
rlabel metal2 s 80044 131200 80100 132000 6 wishbone_out[39]
port 412 nsew signal output
rlabel metal2 s 52628 131200 52684 132000 6 wishbone_out[3]
port 413 nsew signal output
rlabel metal2 s 80872 131200 80928 132000 6 wishbone_out[40]
port 414 nsew signal output
rlabel metal2 s 81608 131200 81664 132000 6 wishbone_out[41]
port 415 nsew signal output
rlabel metal2 s 82344 131200 82400 132000 6 wishbone_out[42]
port 416 nsew signal output
rlabel metal2 s 83172 131200 83228 132000 6 wishbone_out[43]
port 417 nsew signal output
rlabel metal2 s 83908 131200 83964 132000 6 wishbone_out[44]
port 418 nsew signal output
rlabel metal2 s 84644 131200 84700 132000 6 wishbone_out[45]
port 419 nsew signal output
rlabel metal2 s 85472 131200 85528 132000 6 wishbone_out[46]
port 420 nsew signal output
rlabel metal2 s 86208 131200 86264 132000 6 wishbone_out[47]
port 421 nsew signal output
rlabel metal2 s 86944 131200 87000 132000 6 wishbone_out[48]
port 422 nsew signal output
rlabel metal2 s 87680 131200 87736 132000 6 wishbone_out[49]
port 423 nsew signal output
rlabel metal2 s 53364 131200 53420 132000 6 wishbone_out[4]
port 424 nsew signal output
rlabel metal2 s 88508 131200 88564 132000 6 wishbone_out[50]
port 425 nsew signal output
rlabel metal2 s 89244 131200 89300 132000 6 wishbone_out[51]
port 426 nsew signal output
rlabel metal2 s 89980 131200 90036 132000 6 wishbone_out[52]
port 427 nsew signal output
rlabel metal2 s 90808 131200 90864 132000 6 wishbone_out[53]
port 428 nsew signal output
rlabel metal2 s 91544 131200 91600 132000 6 wishbone_out[54]
port 429 nsew signal output
rlabel metal2 s 92280 131200 92336 132000 6 wishbone_out[55]
port 430 nsew signal output
rlabel metal2 s 93016 131200 93072 132000 6 wishbone_out[56]
port 431 nsew signal output
rlabel metal2 s 93844 131200 93900 132000 6 wishbone_out[57]
port 432 nsew signal output
rlabel metal2 s 94580 131200 94636 132000 6 wishbone_out[58]
port 433 nsew signal output
rlabel metal2 s 95316 131200 95372 132000 6 wishbone_out[59]
port 434 nsew signal output
rlabel metal2 s 54100 131200 54156 132000 6 wishbone_out[5]
port 435 nsew signal output
rlabel metal2 s 96144 131200 96200 132000 6 wishbone_out[60]
port 436 nsew signal output
rlabel metal2 s 96880 131200 96936 132000 6 wishbone_out[61]
port 437 nsew signal output
rlabel metal2 s 97616 131200 97672 132000 6 wishbone_out[62]
port 438 nsew signal output
rlabel metal2 s 98444 131200 98500 132000 6 wishbone_out[63]
port 439 nsew signal output
rlabel metal2 s 99180 131200 99236 132000 6 wishbone_out[64]
port 440 nsew signal output
rlabel metal2 s 99916 131200 99972 132000 6 wishbone_out[65]
port 441 nsew signal output
rlabel metal2 s 100652 131200 100708 132000 6 wishbone_out[66]
port 442 nsew signal output
rlabel metal2 s 101480 131200 101536 132000 6 wishbone_out[67]
port 443 nsew signal output
rlabel metal2 s 102216 131200 102272 132000 6 wishbone_out[68]
port 444 nsew signal output
rlabel metal2 s 102952 131200 103008 132000 6 wishbone_out[69]
port 445 nsew signal output
rlabel metal2 s 54928 131200 54984 132000 6 wishbone_out[6]
port 446 nsew signal output
rlabel metal2 s 103780 131200 103836 132000 6 wishbone_out[70]
port 447 nsew signal output
rlabel metal2 s 104516 131200 104572 132000 6 wishbone_out[71]
port 448 nsew signal output
rlabel metal2 s 105252 131200 105308 132000 6 wishbone_out[72]
port 449 nsew signal output
rlabel metal2 s 105988 131200 106044 132000 6 wishbone_out[73]
port 450 nsew signal output
rlabel metal2 s 106816 131200 106872 132000 6 wishbone_out[74]
port 451 nsew signal output
rlabel metal2 s 107552 131200 107608 132000 6 wishbone_out[75]
port 452 nsew signal output
rlabel metal2 s 108288 131200 108344 132000 6 wishbone_out[76]
port 453 nsew signal output
rlabel metal2 s 109116 131200 109172 132000 6 wishbone_out[77]
port 454 nsew signal output
rlabel metal2 s 109852 131200 109908 132000 6 wishbone_out[78]
port 455 nsew signal output
rlabel metal2 s 110588 131200 110644 132000 6 wishbone_out[79]
port 456 nsew signal output
rlabel metal2 s 55664 131200 55720 132000 6 wishbone_out[7]
port 457 nsew signal output
rlabel metal2 s 111416 131200 111472 132000 6 wishbone_out[80]
port 458 nsew signal output
rlabel metal2 s 112152 131200 112208 132000 6 wishbone_out[81]
port 459 nsew signal output
rlabel metal2 s 112888 131200 112944 132000 6 wishbone_out[82]
port 460 nsew signal output
rlabel metal2 s 113624 131200 113680 132000 6 wishbone_out[83]
port 461 nsew signal output
rlabel metal2 s 114452 131200 114508 132000 6 wishbone_out[84]
port 462 nsew signal output
rlabel metal2 s 115188 131200 115244 132000 6 wishbone_out[85]
port 463 nsew signal output
rlabel metal2 s 115924 131200 115980 132000 6 wishbone_out[86]
port 464 nsew signal output
rlabel metal2 s 116752 131200 116808 132000 6 wishbone_out[87]
port 465 nsew signal output
rlabel metal2 s 117488 131200 117544 132000 6 wishbone_out[88]
port 466 nsew signal output
rlabel metal2 s 118224 131200 118280 132000 6 wishbone_out[89]
port 467 nsew signal output
rlabel metal2 s 56400 131200 56456 132000 6 wishbone_out[8]
port 468 nsew signal output
rlabel metal2 s 118960 131200 119016 132000 6 wishbone_out[90]
port 469 nsew signal output
rlabel metal2 s 119788 131200 119844 132000 6 wishbone_out[91]
port 470 nsew signal output
rlabel metal2 s 120524 131200 120580 132000 6 wishbone_out[92]
port 471 nsew signal output
rlabel metal2 s 121260 131200 121316 132000 6 wishbone_out[93]
port 472 nsew signal output
rlabel metal2 s 122088 131200 122144 132000 6 wishbone_out[94]
port 473 nsew signal output
rlabel metal2 s 122824 131200 122880 132000 6 wishbone_out[95]
port 474 nsew signal output
rlabel metal2 s 123560 131200 123616 132000 6 wishbone_out[96]
port 475 nsew signal output
rlabel metal2 s 124388 131200 124444 132000 6 wishbone_out[97]
port 476 nsew signal output
rlabel metal2 s 125124 131200 125180 132000 6 wishbone_out[98]
port 477 nsew signal output
rlabel metal2 s 125860 131200 125916 132000 6 wishbone_out[99]
port 478 nsew signal output
rlabel metal2 s 57228 131200 57284 132000 6 wishbone_out[9]
port 479 nsew signal output
rlabel metal4 s 126706 2128 127026 129520 6 vccd1
port 480 nsew power bidirectional
rlabel metal4 s 95986 2128 96306 129520 6 vccd1
port 481 nsew power bidirectional
rlabel metal4 s 65266 2128 65586 129520 6 vccd1
port 482 nsew power bidirectional
rlabel metal4 s 34546 2128 34866 129520 6 vccd1
port 483 nsew power bidirectional
rlabel metal4 s 3826 2128 4146 129520 6 vccd1
port 484 nsew power bidirectional
rlabel metal4 s 111346 2128 111666 129520 6 vssd1
port 485 nsew ground bidirectional
rlabel metal4 s 80626 2128 80946 129520 6 vssd1
port 486 nsew ground bidirectional
rlabel metal4 s 49906 2128 50226 129520 6 vssd1
port 487 nsew ground bidirectional
rlabel metal4 s 19186 2128 19506 129520 6 vssd1
port 488 nsew ground bidirectional
rlabel metal4 s 127366 2176 127686 129472 6 vccd2
port 489 nsew power bidirectional
rlabel metal4 s 96646 2176 96966 129472 6 vccd2
port 490 nsew power bidirectional
rlabel metal4 s 65926 2176 66246 129472 6 vccd2
port 491 nsew power bidirectional
rlabel metal4 s 35206 2176 35526 129472 6 vccd2
port 492 nsew power bidirectional
rlabel metal4 s 4486 2176 4806 129472 6 vccd2
port 493 nsew power bidirectional
rlabel metal4 s 112006 2176 112326 129472 6 vssd2
port 494 nsew ground bidirectional
rlabel metal4 s 81286 2176 81606 129472 6 vssd2
port 495 nsew ground bidirectional
rlabel metal4 s 50566 2176 50886 129472 6 vssd2
port 496 nsew ground bidirectional
rlabel metal4 s 19846 2176 20166 129472 6 vssd2
port 497 nsew ground bidirectional
rlabel metal4 s 128026 2176 128346 129472 6 vdda1
port 498 nsew power bidirectional
rlabel metal4 s 97306 2176 97626 129472 6 vdda1
port 499 nsew power bidirectional
rlabel metal4 s 66586 2176 66906 129472 6 vdda1
port 500 nsew power bidirectional
rlabel metal4 s 35866 2176 36186 129472 6 vdda1
port 501 nsew power bidirectional
rlabel metal4 s 5146 2176 5466 129472 6 vdda1
port 502 nsew power bidirectional
rlabel metal4 s 112666 2176 112986 129472 6 vssa1
port 503 nsew ground bidirectional
rlabel metal4 s 81946 2176 82266 129472 6 vssa1
port 504 nsew ground bidirectional
rlabel metal4 s 51226 2176 51546 129472 6 vssa1
port 505 nsew ground bidirectional
rlabel metal4 s 20506 2176 20826 129472 6 vssa1
port 506 nsew ground bidirectional
rlabel metal4 s 128686 2176 129006 129472 6 vdda2
port 507 nsew power bidirectional
rlabel metal4 s 97966 2176 98286 129472 6 vdda2
port 508 nsew power bidirectional
rlabel metal4 s 67246 2176 67566 129472 6 vdda2
port 509 nsew power bidirectional
rlabel metal4 s 36526 2176 36846 129472 6 vdda2
port 510 nsew power bidirectional
rlabel metal4 s 5806 2176 6126 129472 6 vdda2
port 511 nsew power bidirectional
rlabel metal4 s 113326 2176 113646 129472 6 vssa2
port 512 nsew ground bidirectional
rlabel metal4 s 82606 2176 82926 129472 6 vssa2
port 513 nsew ground bidirectional
rlabel metal4 s 51886 2176 52206 129472 6 vssa2
port 514 nsew ground bidirectional
rlabel metal4 s 21166 2176 21486 129472 6 vssa2
port 515 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 131618 132000
string LEFview TRUE
<< end >>
