magic
tech sky130A
magscale 1 2
timestamp 1608844419
<< obsli1 >>
rect 1104 791 194856 192313
<< obsm1 >>
rect 1104 760 194856 193784
<< metal2 >>
rect 386 193832 442 194632
rect 1214 193832 1270 194632
rect 2134 193832 2190 194632
rect 3054 193832 3110 194632
rect 3974 193832 4030 194632
rect 4894 193832 4950 194632
rect 5722 193832 5778 194632
rect 6642 193832 6698 194632
rect 7562 193832 7618 194632
rect 8482 193832 8538 194632
rect 9402 193832 9458 194632
rect 10230 193832 10286 194632
rect 11150 193832 11206 194632
rect 12070 193832 12126 194632
rect 12990 193832 13046 194632
rect 13910 193832 13966 194632
rect 14830 193832 14886 194632
rect 15658 193832 15714 194632
rect 16578 193832 16634 194632
rect 17498 193832 17554 194632
rect 18418 193832 18474 194632
rect 19338 193832 19394 194632
rect 20166 193832 20222 194632
rect 21086 193832 21142 194632
rect 22006 193832 22062 194632
rect 22926 193832 22982 194632
rect 23846 193832 23902 194632
rect 24766 193832 24822 194632
rect 25594 193832 25650 194632
rect 26514 193832 26570 194632
rect 27434 193832 27490 194632
rect 28354 193832 28410 194632
rect 29274 193832 29330 194632
rect 30102 193832 30158 194632
rect 31022 193832 31078 194632
rect 31942 193832 31998 194632
rect 32862 193832 32918 194632
rect 33782 193832 33838 194632
rect 34610 193832 34666 194632
rect 35530 193832 35586 194632
rect 36450 193832 36506 194632
rect 37370 193832 37426 194632
rect 38290 193832 38346 194632
rect 39210 193832 39266 194632
rect 40038 193832 40094 194632
rect 40958 193832 41014 194632
rect 41878 193832 41934 194632
rect 42798 193832 42854 194632
rect 43718 193832 43774 194632
rect 44546 193832 44602 194632
rect 45466 193832 45522 194632
rect 46386 193832 46442 194632
rect 47306 193832 47362 194632
rect 48226 193832 48282 194632
rect 49146 193832 49202 194632
rect 49974 193832 50030 194632
rect 50894 193832 50950 194632
rect 51814 193832 51870 194632
rect 52734 193832 52790 194632
rect 53654 193832 53710 194632
rect 54482 193832 54538 194632
rect 55402 193832 55458 194632
rect 56322 193832 56378 194632
rect 57242 193832 57298 194632
rect 58162 193832 58218 194632
rect 59082 193832 59138 194632
rect 59910 193832 59966 194632
rect 60830 193832 60886 194632
rect 61750 193832 61806 194632
rect 62670 193832 62726 194632
rect 63590 193832 63646 194632
rect 64418 193832 64474 194632
rect 65338 193832 65394 194632
rect 66258 193832 66314 194632
rect 67178 193832 67234 194632
rect 68098 193832 68154 194632
rect 68926 193832 68982 194632
rect 69846 193832 69902 194632
rect 70766 193832 70822 194632
rect 71686 193832 71742 194632
rect 72606 193832 72662 194632
rect 73526 193832 73582 194632
rect 74354 193832 74410 194632
rect 75274 193832 75330 194632
rect 76194 193832 76250 194632
rect 77114 193832 77170 194632
rect 78034 193832 78090 194632
rect 78862 193832 78918 194632
rect 79782 193832 79838 194632
rect 80702 193832 80758 194632
rect 81622 193832 81678 194632
rect 82542 193832 82598 194632
rect 83462 193832 83518 194632
rect 84290 193832 84346 194632
rect 85210 193832 85266 194632
rect 86130 193832 86186 194632
rect 87050 193832 87106 194632
rect 87970 193832 88026 194632
rect 88798 193832 88854 194632
rect 89718 193832 89774 194632
rect 90638 193832 90694 194632
rect 91558 193832 91614 194632
rect 92478 193832 92534 194632
rect 93398 193832 93454 194632
rect 94226 193832 94282 194632
rect 95146 193832 95202 194632
rect 96066 193832 96122 194632
rect 96986 193832 97042 194632
rect 97906 193832 97962 194632
rect 98734 193832 98790 194632
rect 99654 193832 99710 194632
rect 100574 193832 100630 194632
rect 101494 193832 101550 194632
rect 102414 193832 102470 194632
rect 103242 193832 103298 194632
rect 104162 193832 104218 194632
rect 105082 193832 105138 194632
rect 106002 193832 106058 194632
rect 106922 193832 106978 194632
rect 107842 193832 107898 194632
rect 108670 193832 108726 194632
rect 109590 193832 109646 194632
rect 110510 193832 110566 194632
rect 111430 193832 111486 194632
rect 112350 193832 112406 194632
rect 113178 193832 113234 194632
rect 114098 193832 114154 194632
rect 115018 193832 115074 194632
rect 115938 193832 115994 194632
rect 116858 193832 116914 194632
rect 117778 193832 117834 194632
rect 118606 193832 118662 194632
rect 119526 193832 119582 194632
rect 120446 193832 120502 194632
rect 121366 193832 121422 194632
rect 122286 193832 122342 194632
rect 123114 193832 123170 194632
rect 124034 193832 124090 194632
rect 124954 193832 125010 194632
rect 125874 193832 125930 194632
rect 126794 193832 126850 194632
rect 127714 193832 127770 194632
rect 128542 193832 128598 194632
rect 129462 193832 129518 194632
rect 130382 193832 130438 194632
rect 131302 193832 131358 194632
rect 132222 193832 132278 194632
rect 133050 193832 133106 194632
rect 133970 193832 134026 194632
rect 134890 193832 134946 194632
rect 135810 193832 135866 194632
rect 136730 193832 136786 194632
rect 137558 193832 137614 194632
rect 138478 193832 138534 194632
rect 139398 193832 139454 194632
rect 140318 193832 140374 194632
rect 141238 193832 141294 194632
rect 142158 193832 142214 194632
rect 142986 193832 143042 194632
rect 143906 193832 143962 194632
rect 144826 193832 144882 194632
rect 145746 193832 145802 194632
rect 146666 193832 146722 194632
rect 147494 193832 147550 194632
rect 148414 193832 148470 194632
rect 149334 193832 149390 194632
rect 150254 193832 150310 194632
rect 151174 193832 151230 194632
rect 152094 193832 152150 194632
rect 152922 193832 152978 194632
rect 153842 193832 153898 194632
rect 154762 193832 154818 194632
rect 155682 193832 155738 194632
rect 156602 193832 156658 194632
rect 157430 193832 157486 194632
rect 158350 193832 158406 194632
rect 159270 193832 159326 194632
rect 160190 193832 160246 194632
rect 161110 193832 161166 194632
rect 162030 193832 162086 194632
rect 162858 193832 162914 194632
rect 163778 193832 163834 194632
rect 164698 193832 164754 194632
rect 165618 193832 165674 194632
rect 166538 193832 166594 194632
rect 167366 193832 167422 194632
rect 168286 193832 168342 194632
rect 169206 193832 169262 194632
rect 170126 193832 170182 194632
rect 171046 193832 171102 194632
rect 171874 193832 171930 194632
rect 172794 193832 172850 194632
rect 173714 193832 173770 194632
rect 174634 193832 174690 194632
rect 175554 193832 175610 194632
rect 176474 193832 176530 194632
rect 177302 193832 177358 194632
rect 178222 193832 178278 194632
rect 179142 193832 179198 194632
rect 180062 193832 180118 194632
rect 180982 193832 181038 194632
rect 181810 193832 181866 194632
rect 182730 193832 182786 194632
rect 183650 193832 183706 194632
rect 184570 193832 184626 194632
rect 185490 193832 185546 194632
rect 186410 193832 186466 194632
rect 187238 193832 187294 194632
rect 188158 193832 188214 194632
rect 189078 193832 189134 194632
rect 189998 193832 190054 194632
rect 190918 193832 190974 194632
rect 191746 193832 191802 194632
rect 192666 193832 192722 194632
rect 193586 193832 193642 194632
rect 194506 193832 194562 194632
rect 195426 193832 195482 194632
<< obsm2 >>
rect 498 193776 1158 193832
rect 1326 193776 2078 193832
rect 2246 193776 2998 193832
rect 3166 193776 3918 193832
rect 4086 193776 4838 193832
rect 5006 193776 5666 193832
rect 5834 193776 6586 193832
rect 6754 193776 7506 193832
rect 7674 193776 8426 193832
rect 8594 193776 9346 193832
rect 9514 193776 10174 193832
rect 10342 193776 11094 193832
rect 11262 193776 12014 193832
rect 12182 193776 12934 193832
rect 13102 193776 13854 193832
rect 14022 193776 14774 193832
rect 14942 193776 15602 193832
rect 15770 193776 16522 193832
rect 16690 193776 17442 193832
rect 17610 193776 18362 193832
rect 18530 193776 19282 193832
rect 19450 193776 20110 193832
rect 20278 193776 21030 193832
rect 21198 193776 21950 193832
rect 22118 193776 22870 193832
rect 23038 193776 23790 193832
rect 23958 193776 24710 193832
rect 24878 193776 25538 193832
rect 25706 193776 26458 193832
rect 26626 193776 27378 193832
rect 27546 193776 28298 193832
rect 28466 193776 29218 193832
rect 29386 193776 30046 193832
rect 30214 193776 30966 193832
rect 31134 193776 31886 193832
rect 32054 193776 32806 193832
rect 32974 193776 33726 193832
rect 33894 193776 34554 193832
rect 34722 193776 35474 193832
rect 35642 193776 36394 193832
rect 36562 193776 37314 193832
rect 37482 193776 38234 193832
rect 38402 193776 39154 193832
rect 39322 193776 39982 193832
rect 40150 193776 40902 193832
rect 41070 193776 41822 193832
rect 41990 193776 42742 193832
rect 42910 193776 43662 193832
rect 43830 193776 44490 193832
rect 44658 193776 45410 193832
rect 45578 193776 46330 193832
rect 46498 193776 47250 193832
rect 47418 193776 48170 193832
rect 48338 193776 49090 193832
rect 49258 193776 49918 193832
rect 50086 193776 50838 193832
rect 51006 193776 51758 193832
rect 51926 193776 52678 193832
rect 52846 193776 53598 193832
rect 53766 193776 54426 193832
rect 54594 193776 55346 193832
rect 55514 193776 56266 193832
rect 56434 193776 57186 193832
rect 57354 193776 58106 193832
rect 58274 193776 59026 193832
rect 59194 193776 59854 193832
rect 60022 193776 60774 193832
rect 60942 193776 61694 193832
rect 61862 193776 62614 193832
rect 62782 193776 63534 193832
rect 63702 193776 64362 193832
rect 64530 193776 65282 193832
rect 65450 193776 66202 193832
rect 66370 193776 67122 193832
rect 67290 193776 68042 193832
rect 68210 193776 68870 193832
rect 69038 193776 69790 193832
rect 69958 193776 70710 193832
rect 70878 193776 71630 193832
rect 71798 193776 72550 193832
rect 72718 193776 73470 193832
rect 73638 193776 74298 193832
rect 74466 193776 75218 193832
rect 75386 193776 76138 193832
rect 76306 193776 77058 193832
rect 77226 193776 77978 193832
rect 78146 193776 78806 193832
rect 78974 193776 79726 193832
rect 79894 193776 80646 193832
rect 80814 193776 81566 193832
rect 81734 193776 82486 193832
rect 82654 193776 83406 193832
rect 83574 193776 84234 193832
rect 84402 193776 85154 193832
rect 85322 193776 86074 193832
rect 86242 193776 86994 193832
rect 87162 193776 87914 193832
rect 88082 193776 88742 193832
rect 88910 193776 89662 193832
rect 89830 193776 90582 193832
rect 90750 193776 91502 193832
rect 91670 193776 92422 193832
rect 92590 193776 93342 193832
rect 93510 193776 94170 193832
rect 94338 193776 95090 193832
rect 95258 193776 96010 193832
rect 96178 193776 96930 193832
rect 97098 193776 97850 193832
rect 98018 193776 98678 193832
rect 98846 193776 99598 193832
rect 99766 193776 100518 193832
rect 100686 193776 101438 193832
rect 101606 193776 102358 193832
rect 102526 193776 103186 193832
rect 103354 193776 104106 193832
rect 104274 193776 105026 193832
rect 105194 193776 105946 193832
rect 106114 193776 106866 193832
rect 107034 193776 107786 193832
rect 107954 193776 108614 193832
rect 108782 193776 109534 193832
rect 109702 193776 110454 193832
rect 110622 193776 111374 193832
rect 111542 193776 112294 193832
rect 112462 193776 113122 193832
rect 113290 193776 114042 193832
rect 114210 193776 114962 193832
rect 115130 193776 115882 193832
rect 116050 193776 116802 193832
rect 116970 193776 117722 193832
rect 117890 193776 118550 193832
rect 118718 193776 119470 193832
rect 119638 193776 120390 193832
rect 120558 193776 121310 193832
rect 121478 193776 122230 193832
rect 122398 193776 123058 193832
rect 123226 193776 123978 193832
rect 124146 193776 124898 193832
rect 125066 193776 125818 193832
rect 125986 193776 126738 193832
rect 126906 193776 127658 193832
rect 127826 193776 128486 193832
rect 128654 193776 129406 193832
rect 129574 193776 130326 193832
rect 130494 193776 131246 193832
rect 131414 193776 132166 193832
rect 132334 193776 132994 193832
rect 133162 193776 133914 193832
rect 134082 193776 134834 193832
rect 135002 193776 135754 193832
rect 135922 193776 136674 193832
rect 136842 193776 137502 193832
rect 137670 193776 138422 193832
rect 138590 193776 139342 193832
rect 139510 193776 140262 193832
rect 140430 193776 141182 193832
rect 141350 193776 142102 193832
rect 142270 193776 142930 193832
rect 143098 193776 143850 193832
rect 144018 193776 144770 193832
rect 144938 193776 145690 193832
rect 145858 193776 146610 193832
rect 146778 193776 147438 193832
rect 147606 193776 148358 193832
rect 148526 193776 149278 193832
rect 149446 193776 150198 193832
rect 150366 193776 151118 193832
rect 151286 193776 152038 193832
rect 152206 193776 152866 193832
rect 153034 193776 153786 193832
rect 153954 193776 154706 193832
rect 154874 193776 155626 193832
rect 155794 193776 156546 193832
rect 156714 193776 157374 193832
rect 157542 193776 158294 193832
rect 158462 193776 159214 193832
rect 159382 193776 160134 193832
rect 160302 193776 161054 193832
rect 161222 193776 161974 193832
rect 162142 193776 162802 193832
rect 162970 193776 163722 193832
rect 163890 193776 164642 193832
rect 164810 193776 165562 193832
rect 165730 193776 166482 193832
rect 166650 193776 167310 193832
rect 167478 193776 168230 193832
rect 168398 193776 169150 193832
rect 169318 193776 170070 193832
rect 170238 193776 170990 193832
rect 171158 193776 171818 193832
rect 171986 193776 172738 193832
rect 172906 193776 173658 193832
rect 173826 193776 174578 193832
rect 174746 193776 175498 193832
rect 175666 193776 176418 193832
rect 176586 193776 177246 193832
rect 177414 193776 178166 193832
rect 178334 193776 179086 193832
rect 179254 193776 180006 193832
rect 180174 193776 180926 193832
rect 181094 193776 181754 193832
rect 181922 193776 182674 193832
rect 182842 193776 183594 193832
rect 183762 193776 184514 193832
rect 184682 193776 185434 193832
rect 185602 193776 186354 193832
rect 186522 193776 187182 193832
rect 187350 193776 188102 193832
rect 188270 193776 189022 193832
rect 189190 193776 189942 193832
rect 190110 193776 190862 193832
rect 191030 193776 191690 193832
rect 191858 193776 192610 193832
rect 192778 193776 193530 193832
rect 193698 193776 194450 193832
rect 194618 193776 195370 193832
rect 386 760 195468 193776
<< metal3 >>
rect 0 193120 800 193240
rect 0 190400 800 190520
rect 0 187680 800 187800
rect 0 184960 800 185080
rect 0 182240 800 182360
rect 0 179520 800 179640
rect 0 176800 800 176920
rect 0 174080 800 174200
rect 0 171360 800 171480
rect 0 168640 800 168760
rect 0 165920 800 166040
rect 0 163200 800 163320
rect 0 160480 800 160600
rect 0 157760 800 157880
rect 0 155040 800 155160
rect 0 152320 800 152440
rect 0 149600 800 149720
rect 0 146880 800 147000
rect 0 144160 800 144280
rect 0 141440 800 141560
rect 0 138720 800 138840
rect 0 136000 800 136120
rect 0 133280 800 133400
rect 0 130560 800 130680
rect 0 127840 800 127960
rect 0 125120 800 125240
rect 0 122400 800 122520
rect 0 119680 800 119800
rect 0 116960 800 117080
rect 0 114240 800 114360
rect 0 111520 800 111640
rect 0 108800 800 108920
rect 0 106080 800 106200
rect 0 103360 800 103480
rect 0 100640 800 100760
rect 0 97920 800 98040
rect 0 95200 800 95320
rect 0 92480 800 92600
rect 0 89760 800 89880
rect 0 87040 800 87160
rect 0 84320 800 84440
rect 0 81600 800 81720
rect 0 78880 800 79000
rect 0 76160 800 76280
rect 0 73440 800 73560
rect 0 70720 800 70840
rect 0 68000 800 68120
rect 0 65280 800 65400
rect 0 62560 800 62680
rect 0 59840 800 59960
rect 0 57120 800 57240
rect 0 54400 800 54520
rect 0 51680 800 51800
rect 0 48960 800 49080
rect 0 46240 800 46360
rect 0 43520 800 43640
rect 0 40800 800 40920
rect 0 38080 800 38200
rect 0 35360 800 35480
rect 0 32640 800 32760
rect 0 29920 800 30040
rect 0 27200 800 27320
rect 0 24480 800 24600
rect 0 21760 800 21880
rect 0 19040 800 19160
rect 0 16320 800 16440
rect 0 13600 800 13720
rect 0 10880 800 11000
rect 0 8160 800 8280
rect 0 5440 800 5560
rect 0 2720 800 2840
rect 0 0 800 120
<< obsm3 >>
rect 880 193040 194659 193213
rect 381 190600 194659 193040
rect 880 190320 194659 190600
rect 381 187880 194659 190320
rect 880 187600 194659 187880
rect 381 185160 194659 187600
rect 880 184880 194659 185160
rect 381 182440 194659 184880
rect 880 182160 194659 182440
rect 381 179720 194659 182160
rect 880 179440 194659 179720
rect 381 177000 194659 179440
rect 880 176720 194659 177000
rect 381 174280 194659 176720
rect 880 174000 194659 174280
rect 381 171560 194659 174000
rect 880 171280 194659 171560
rect 381 168840 194659 171280
rect 880 168560 194659 168840
rect 381 166120 194659 168560
rect 880 165840 194659 166120
rect 381 163400 194659 165840
rect 880 163120 194659 163400
rect 381 160680 194659 163120
rect 880 160400 194659 160680
rect 381 157960 194659 160400
rect 880 157680 194659 157960
rect 381 155240 194659 157680
rect 880 154960 194659 155240
rect 381 152520 194659 154960
rect 880 152240 194659 152520
rect 381 149800 194659 152240
rect 880 149520 194659 149800
rect 381 147080 194659 149520
rect 880 146800 194659 147080
rect 381 144360 194659 146800
rect 880 144080 194659 144360
rect 381 141640 194659 144080
rect 880 141360 194659 141640
rect 381 138920 194659 141360
rect 880 138640 194659 138920
rect 381 136200 194659 138640
rect 880 135920 194659 136200
rect 381 133480 194659 135920
rect 880 133200 194659 133480
rect 381 130760 194659 133200
rect 880 130480 194659 130760
rect 381 128040 194659 130480
rect 880 127760 194659 128040
rect 381 125320 194659 127760
rect 880 125040 194659 125320
rect 381 122600 194659 125040
rect 880 122320 194659 122600
rect 381 119880 194659 122320
rect 880 119600 194659 119880
rect 381 117160 194659 119600
rect 880 116880 194659 117160
rect 381 114440 194659 116880
rect 880 114160 194659 114440
rect 381 111720 194659 114160
rect 880 111440 194659 111720
rect 381 109000 194659 111440
rect 880 108720 194659 109000
rect 381 106280 194659 108720
rect 880 106000 194659 106280
rect 381 103560 194659 106000
rect 880 103280 194659 103560
rect 381 100840 194659 103280
rect 880 100560 194659 100840
rect 381 98120 194659 100560
rect 880 97840 194659 98120
rect 381 95400 194659 97840
rect 880 95120 194659 95400
rect 381 92680 194659 95120
rect 880 92400 194659 92680
rect 381 89960 194659 92400
rect 880 89680 194659 89960
rect 381 87240 194659 89680
rect 880 86960 194659 87240
rect 381 84520 194659 86960
rect 880 84240 194659 84520
rect 381 81800 194659 84240
rect 880 81520 194659 81800
rect 381 79080 194659 81520
rect 880 78800 194659 79080
rect 381 76360 194659 78800
rect 880 76080 194659 76360
rect 381 73640 194659 76080
rect 880 73360 194659 73640
rect 381 70920 194659 73360
rect 880 70640 194659 70920
rect 381 68200 194659 70640
rect 880 67920 194659 68200
rect 381 65480 194659 67920
rect 880 65200 194659 65480
rect 381 62760 194659 65200
rect 880 62480 194659 62760
rect 381 60040 194659 62480
rect 880 59760 194659 60040
rect 381 57320 194659 59760
rect 880 57040 194659 57320
rect 381 54600 194659 57040
rect 880 54320 194659 54600
rect 381 51880 194659 54320
rect 880 51600 194659 51880
rect 381 49160 194659 51600
rect 880 48880 194659 49160
rect 381 46440 194659 48880
rect 880 46160 194659 46440
rect 381 43720 194659 46160
rect 880 43440 194659 43720
rect 381 41000 194659 43440
rect 880 40720 194659 41000
rect 381 38280 194659 40720
rect 880 38000 194659 38280
rect 381 35560 194659 38000
rect 880 35280 194659 35560
rect 381 32840 194659 35280
rect 880 32560 194659 32840
rect 381 30120 194659 32560
rect 880 29840 194659 30120
rect 381 27400 194659 29840
rect 880 27120 194659 27400
rect 381 24680 194659 27120
rect 880 24400 194659 24680
rect 381 21960 194659 24400
rect 880 21680 194659 21960
rect 381 19240 194659 21680
rect 880 18960 194659 19240
rect 381 16520 194659 18960
rect 880 16240 194659 16520
rect 381 13800 194659 16240
rect 880 13520 194659 13800
rect 381 11080 194659 13520
rect 880 10800 194659 11080
rect 381 8360 194659 10800
rect 880 8080 194659 8360
rect 381 5640 194659 8080
rect 880 5360 194659 5640
rect 381 2920 194659 5360
rect 880 2640 194659 2920
rect 381 200 194659 2640
rect 880 28 194659 200
<< metal4 >>
rect 4208 760 4528 192344
rect 4868 808 5188 192296
rect 5528 808 5848 192296
rect 6188 808 6508 192296
rect 19568 760 19888 192344
rect 20228 808 20548 192296
rect 20888 808 21208 192296
rect 21548 808 21868 192296
rect 34928 760 35248 192344
rect 35588 808 35908 192296
rect 36248 808 36568 192296
rect 36908 808 37228 192296
rect 50288 760 50608 192344
rect 50948 808 51268 192296
rect 51608 808 51928 192296
rect 52268 808 52588 192296
rect 65648 760 65968 192344
rect 66308 808 66628 192296
rect 66968 808 67288 192296
rect 67628 808 67948 192296
rect 81008 760 81328 192344
rect 81668 808 81988 192296
rect 82328 808 82648 192296
rect 82988 808 83308 192296
rect 96368 760 96688 192344
rect 97028 808 97348 192296
rect 97688 808 98008 192296
rect 98348 808 98668 192296
rect 111728 760 112048 192344
rect 112388 808 112708 192296
rect 113048 808 113368 192296
rect 113708 808 114028 192296
rect 127088 760 127408 192344
rect 127748 808 128068 192296
rect 128408 808 128728 192296
rect 129068 808 129388 192296
rect 142448 760 142768 192344
rect 143108 808 143428 192296
rect 143768 808 144088 192296
rect 144428 808 144748 192296
rect 157808 760 158128 192344
rect 158468 808 158788 192296
rect 159128 808 159448 192296
rect 159788 808 160108 192296
rect 173168 760 173488 192344
rect 173828 808 174148 192296
rect 174488 808 174808 192296
rect 175148 808 175468 192296
rect 188528 760 188848 192344
rect 189188 808 189508 192296
rect 189848 808 190168 192296
rect 190508 808 190828 192296
<< obsm4 >>
rect 1715 680 4128 192397
rect 4608 192376 19488 192397
rect 4608 728 4788 192376
rect 5268 728 5448 192376
rect 5928 728 6108 192376
rect 6588 728 19488 192376
rect 19968 192376 34848 192397
rect 4608 680 19488 728
rect 19968 728 20148 192376
rect 20628 728 20808 192376
rect 21288 728 21468 192376
rect 21948 728 34848 192376
rect 35328 192376 50208 192397
rect 19968 680 34848 728
rect 35328 728 35508 192376
rect 35988 728 36168 192376
rect 36648 728 36828 192376
rect 37308 728 50208 192376
rect 50688 192376 65568 192397
rect 35328 680 50208 728
rect 50688 728 50868 192376
rect 51348 728 51528 192376
rect 52008 728 52188 192376
rect 52668 728 65568 192376
rect 66048 192376 80928 192397
rect 50688 680 65568 728
rect 66048 728 66228 192376
rect 66708 728 66888 192376
rect 67368 728 67548 192376
rect 68028 728 80928 192376
rect 81408 192376 96288 192397
rect 66048 680 80928 728
rect 81408 728 81588 192376
rect 82068 728 82248 192376
rect 82728 728 82908 192376
rect 83388 728 96288 192376
rect 96768 192376 111648 192397
rect 81408 680 96288 728
rect 96768 728 96948 192376
rect 97428 728 97608 192376
rect 98088 728 98268 192376
rect 98748 728 111648 192376
rect 112128 192376 127008 192397
rect 96768 680 111648 728
rect 112128 728 112308 192376
rect 112788 728 112968 192376
rect 113448 728 113628 192376
rect 114108 728 127008 192376
rect 127488 192376 142368 192397
rect 112128 680 127008 728
rect 127488 728 127668 192376
rect 128148 728 128328 192376
rect 128808 728 128988 192376
rect 129468 728 142368 192376
rect 142848 192376 157728 192397
rect 127488 680 142368 728
rect 142848 728 143028 192376
rect 143508 728 143688 192376
rect 144168 728 144348 192376
rect 144828 728 157728 192376
rect 158208 192376 173088 192397
rect 142848 680 157728 728
rect 158208 728 158388 192376
rect 158868 728 159048 192376
rect 159528 728 159708 192376
rect 160188 728 173088 192376
rect 173568 192376 188448 192397
rect 158208 680 173088 728
rect 173568 728 173748 192376
rect 174228 728 174408 192376
rect 174888 728 175068 192376
rect 175548 728 188448 192376
rect 188928 192376 192957 192397
rect 173568 680 188448 728
rect 188928 728 189108 192376
rect 189588 728 189768 192376
rect 190248 728 190428 192376
rect 190908 728 192957 192376
rect 188928 680 192957 728
rect 1715 27 192957 680
<< obsm5 >>
rect 71324 110332 73116 110652
<< labels >>
rlabel metal2 s 386 193832 442 194632 6 clk
port 1 nsew signal input
rlabel metal2 s 1214 193832 1270 194632 6 d_in[0]
port 2 nsew signal input
rlabel metal2 s 10230 193832 10286 194632 6 d_in[10]
port 3 nsew signal input
rlabel metal2 s 11150 193832 11206 194632 6 d_in[11]
port 4 nsew signal input
rlabel metal2 s 12070 193832 12126 194632 6 d_in[12]
port 5 nsew signal input
rlabel metal2 s 12990 193832 13046 194632 6 d_in[13]
port 6 nsew signal input
rlabel metal2 s 13910 193832 13966 194632 6 d_in[14]
port 7 nsew signal input
rlabel metal2 s 14830 193832 14886 194632 6 d_in[15]
port 8 nsew signal input
rlabel metal2 s 15658 193832 15714 194632 6 d_in[16]
port 9 nsew signal input
rlabel metal2 s 16578 193832 16634 194632 6 d_in[17]
port 10 nsew signal input
rlabel metal2 s 17498 193832 17554 194632 6 d_in[18]
port 11 nsew signal input
rlabel metal2 s 18418 193832 18474 194632 6 d_in[19]
port 12 nsew signal input
rlabel metal2 s 2134 193832 2190 194632 6 d_in[1]
port 13 nsew signal input
rlabel metal2 s 19338 193832 19394 194632 6 d_in[20]
port 14 nsew signal input
rlabel metal2 s 20166 193832 20222 194632 6 d_in[21]
port 15 nsew signal input
rlabel metal2 s 21086 193832 21142 194632 6 d_in[22]
port 16 nsew signal input
rlabel metal2 s 22006 193832 22062 194632 6 d_in[23]
port 17 nsew signal input
rlabel metal2 s 3054 193832 3110 194632 6 d_in[2]
port 18 nsew signal input
rlabel metal2 s 3974 193832 4030 194632 6 d_in[3]
port 19 nsew signal input
rlabel metal2 s 4894 193832 4950 194632 6 d_in[4]
port 20 nsew signal input
rlabel metal2 s 5722 193832 5778 194632 6 d_in[5]
port 21 nsew signal input
rlabel metal2 s 6642 193832 6698 194632 6 d_in[6]
port 22 nsew signal input
rlabel metal2 s 7562 193832 7618 194632 6 d_in[7]
port 23 nsew signal input
rlabel metal2 s 8482 193832 8538 194632 6 d_in[8]
port 24 nsew signal input
rlabel metal2 s 9402 193832 9458 194632 6 d_in[9]
port 25 nsew signal input
rlabel metal2 s 22926 193832 22982 194632 6 d_out[0]
port 26 nsew signal output
rlabel metal2 s 113178 193832 113234 194632 6 d_out[100]
port 27 nsew signal output
rlabel metal2 s 114098 193832 114154 194632 6 d_out[101]
port 28 nsew signal output
rlabel metal2 s 115018 193832 115074 194632 6 d_out[102]
port 29 nsew signal output
rlabel metal2 s 115938 193832 115994 194632 6 d_out[103]
port 30 nsew signal output
rlabel metal2 s 116858 193832 116914 194632 6 d_out[104]
port 31 nsew signal output
rlabel metal2 s 117778 193832 117834 194632 6 d_out[105]
port 32 nsew signal output
rlabel metal2 s 118606 193832 118662 194632 6 d_out[106]
port 33 nsew signal output
rlabel metal2 s 119526 193832 119582 194632 6 d_out[107]
port 34 nsew signal output
rlabel metal2 s 120446 193832 120502 194632 6 d_out[108]
port 35 nsew signal output
rlabel metal2 s 121366 193832 121422 194632 6 d_out[109]
port 36 nsew signal output
rlabel metal2 s 31942 193832 31998 194632 6 d_out[10]
port 37 nsew signal output
rlabel metal2 s 122286 193832 122342 194632 6 d_out[110]
port 38 nsew signal output
rlabel metal2 s 123114 193832 123170 194632 6 d_out[111]
port 39 nsew signal output
rlabel metal2 s 124034 193832 124090 194632 6 d_out[112]
port 40 nsew signal output
rlabel metal2 s 124954 193832 125010 194632 6 d_out[113]
port 41 nsew signal output
rlabel metal2 s 125874 193832 125930 194632 6 d_out[114]
port 42 nsew signal output
rlabel metal2 s 126794 193832 126850 194632 6 d_out[115]
port 43 nsew signal output
rlabel metal2 s 127714 193832 127770 194632 6 d_out[116]
port 44 nsew signal output
rlabel metal2 s 128542 193832 128598 194632 6 d_out[117]
port 45 nsew signal output
rlabel metal2 s 129462 193832 129518 194632 6 d_out[118]
port 46 nsew signal output
rlabel metal2 s 130382 193832 130438 194632 6 d_out[119]
port 47 nsew signal output
rlabel metal2 s 32862 193832 32918 194632 6 d_out[11]
port 48 nsew signal output
rlabel metal2 s 131302 193832 131358 194632 6 d_out[120]
port 49 nsew signal output
rlabel metal2 s 132222 193832 132278 194632 6 d_out[121]
port 50 nsew signal output
rlabel metal2 s 133050 193832 133106 194632 6 d_out[122]
port 51 nsew signal output
rlabel metal2 s 133970 193832 134026 194632 6 d_out[123]
port 52 nsew signal output
rlabel metal2 s 134890 193832 134946 194632 6 d_out[124]
port 53 nsew signal output
rlabel metal2 s 135810 193832 135866 194632 6 d_out[125]
port 54 nsew signal output
rlabel metal2 s 136730 193832 136786 194632 6 d_out[126]
port 55 nsew signal output
rlabel metal2 s 137558 193832 137614 194632 6 d_out[127]
port 56 nsew signal output
rlabel metal2 s 138478 193832 138534 194632 6 d_out[128]
port 57 nsew signal output
rlabel metal2 s 139398 193832 139454 194632 6 d_out[129]
port 58 nsew signal output
rlabel metal2 s 33782 193832 33838 194632 6 d_out[12]
port 59 nsew signal output
rlabel metal2 s 140318 193832 140374 194632 6 d_out[130]
port 60 nsew signal output
rlabel metal2 s 141238 193832 141294 194632 6 d_out[131]
port 61 nsew signal output
rlabel metal2 s 142158 193832 142214 194632 6 d_out[132]
port 62 nsew signal output
rlabel metal2 s 142986 193832 143042 194632 6 d_out[133]
port 63 nsew signal output
rlabel metal2 s 143906 193832 143962 194632 6 d_out[134]
port 64 nsew signal output
rlabel metal2 s 144826 193832 144882 194632 6 d_out[135]
port 65 nsew signal output
rlabel metal2 s 145746 193832 145802 194632 6 d_out[136]
port 66 nsew signal output
rlabel metal2 s 146666 193832 146722 194632 6 d_out[137]
port 67 nsew signal output
rlabel metal2 s 147494 193832 147550 194632 6 d_out[138]
port 68 nsew signal output
rlabel metal2 s 148414 193832 148470 194632 6 d_out[139]
port 69 nsew signal output
rlabel metal2 s 34610 193832 34666 194632 6 d_out[13]
port 70 nsew signal output
rlabel metal2 s 149334 193832 149390 194632 6 d_out[140]
port 71 nsew signal output
rlabel metal2 s 150254 193832 150310 194632 6 d_out[141]
port 72 nsew signal output
rlabel metal2 s 151174 193832 151230 194632 6 d_out[142]
port 73 nsew signal output
rlabel metal2 s 152094 193832 152150 194632 6 d_out[143]
port 74 nsew signal output
rlabel metal2 s 152922 193832 152978 194632 6 d_out[144]
port 75 nsew signal output
rlabel metal2 s 153842 193832 153898 194632 6 d_out[145]
port 76 nsew signal output
rlabel metal2 s 154762 193832 154818 194632 6 d_out[146]
port 77 nsew signal output
rlabel metal2 s 155682 193832 155738 194632 6 d_out[147]
port 78 nsew signal output
rlabel metal2 s 156602 193832 156658 194632 6 d_out[148]
port 79 nsew signal output
rlabel metal2 s 157430 193832 157486 194632 6 d_out[149]
port 80 nsew signal output
rlabel metal2 s 35530 193832 35586 194632 6 d_out[14]
port 81 nsew signal output
rlabel metal2 s 158350 193832 158406 194632 6 d_out[150]
port 82 nsew signal output
rlabel metal2 s 159270 193832 159326 194632 6 d_out[151]
port 83 nsew signal output
rlabel metal2 s 160190 193832 160246 194632 6 d_out[152]
port 84 nsew signal output
rlabel metal2 s 161110 193832 161166 194632 6 d_out[153]
port 85 nsew signal output
rlabel metal2 s 162030 193832 162086 194632 6 d_out[154]
port 86 nsew signal output
rlabel metal2 s 162858 193832 162914 194632 6 d_out[155]
port 87 nsew signal output
rlabel metal2 s 163778 193832 163834 194632 6 d_out[156]
port 88 nsew signal output
rlabel metal2 s 164698 193832 164754 194632 6 d_out[157]
port 89 nsew signal output
rlabel metal2 s 165618 193832 165674 194632 6 d_out[158]
port 90 nsew signal output
rlabel metal2 s 166538 193832 166594 194632 6 d_out[159]
port 91 nsew signal output
rlabel metal2 s 36450 193832 36506 194632 6 d_out[15]
port 92 nsew signal output
rlabel metal2 s 167366 193832 167422 194632 6 d_out[160]
port 93 nsew signal output
rlabel metal2 s 168286 193832 168342 194632 6 d_out[161]
port 94 nsew signal output
rlabel metal2 s 169206 193832 169262 194632 6 d_out[162]
port 95 nsew signal output
rlabel metal2 s 170126 193832 170182 194632 6 d_out[163]
port 96 nsew signal output
rlabel metal2 s 171046 193832 171102 194632 6 d_out[164]
port 97 nsew signal output
rlabel metal2 s 171874 193832 171930 194632 6 d_out[165]
port 98 nsew signal output
rlabel metal2 s 172794 193832 172850 194632 6 d_out[166]
port 99 nsew signal output
rlabel metal2 s 173714 193832 173770 194632 6 d_out[167]
port 100 nsew signal output
rlabel metal2 s 174634 193832 174690 194632 6 d_out[168]
port 101 nsew signal output
rlabel metal2 s 175554 193832 175610 194632 6 d_out[169]
port 102 nsew signal output
rlabel metal2 s 37370 193832 37426 194632 6 d_out[16]
port 103 nsew signal output
rlabel metal2 s 176474 193832 176530 194632 6 d_out[170]
port 104 nsew signal output
rlabel metal2 s 177302 193832 177358 194632 6 d_out[171]
port 105 nsew signal output
rlabel metal2 s 178222 193832 178278 194632 6 d_out[172]
port 106 nsew signal output
rlabel metal2 s 179142 193832 179198 194632 6 d_out[173]
port 107 nsew signal output
rlabel metal2 s 180062 193832 180118 194632 6 d_out[174]
port 108 nsew signal output
rlabel metal2 s 180982 193832 181038 194632 6 d_out[175]
port 109 nsew signal output
rlabel metal2 s 181810 193832 181866 194632 6 d_out[176]
port 110 nsew signal output
rlabel metal2 s 182730 193832 182786 194632 6 d_out[177]
port 111 nsew signal output
rlabel metal2 s 183650 193832 183706 194632 6 d_out[178]
port 112 nsew signal output
rlabel metal2 s 184570 193832 184626 194632 6 d_out[179]
port 113 nsew signal output
rlabel metal2 s 38290 193832 38346 194632 6 d_out[17]
port 114 nsew signal output
rlabel metal2 s 185490 193832 185546 194632 6 d_out[180]
port 115 nsew signal output
rlabel metal2 s 186410 193832 186466 194632 6 d_out[181]
port 116 nsew signal output
rlabel metal2 s 187238 193832 187294 194632 6 d_out[182]
port 117 nsew signal output
rlabel metal2 s 188158 193832 188214 194632 6 d_out[183]
port 118 nsew signal output
rlabel metal2 s 189078 193832 189134 194632 6 d_out[184]
port 119 nsew signal output
rlabel metal2 s 189998 193832 190054 194632 6 d_out[185]
port 120 nsew signal output
rlabel metal2 s 190918 193832 190974 194632 6 d_out[186]
port 121 nsew signal output
rlabel metal2 s 191746 193832 191802 194632 6 d_out[187]
port 122 nsew signal output
rlabel metal2 s 192666 193832 192722 194632 6 d_out[188]
port 123 nsew signal output
rlabel metal2 s 193586 193832 193642 194632 6 d_out[189]
port 124 nsew signal output
rlabel metal2 s 39210 193832 39266 194632 6 d_out[18]
port 125 nsew signal output
rlabel metal2 s 194506 193832 194562 194632 6 d_out[190]
port 126 nsew signal output
rlabel metal2 s 195426 193832 195482 194632 6 d_out[191]
port 127 nsew signal output
rlabel metal2 s 40038 193832 40094 194632 6 d_out[19]
port 128 nsew signal output
rlabel metal2 s 23846 193832 23902 194632 6 d_out[1]
port 129 nsew signal output
rlabel metal2 s 40958 193832 41014 194632 6 d_out[20]
port 130 nsew signal output
rlabel metal2 s 41878 193832 41934 194632 6 d_out[21]
port 131 nsew signal output
rlabel metal2 s 42798 193832 42854 194632 6 d_out[22]
port 132 nsew signal output
rlabel metal2 s 43718 193832 43774 194632 6 d_out[23]
port 133 nsew signal output
rlabel metal2 s 44546 193832 44602 194632 6 d_out[24]
port 134 nsew signal output
rlabel metal2 s 45466 193832 45522 194632 6 d_out[25]
port 135 nsew signal output
rlabel metal2 s 46386 193832 46442 194632 6 d_out[26]
port 136 nsew signal output
rlabel metal2 s 47306 193832 47362 194632 6 d_out[27]
port 137 nsew signal output
rlabel metal2 s 48226 193832 48282 194632 6 d_out[28]
port 138 nsew signal output
rlabel metal2 s 49146 193832 49202 194632 6 d_out[29]
port 139 nsew signal output
rlabel metal2 s 24766 193832 24822 194632 6 d_out[2]
port 140 nsew signal output
rlabel metal2 s 49974 193832 50030 194632 6 d_out[30]
port 141 nsew signal output
rlabel metal2 s 50894 193832 50950 194632 6 d_out[31]
port 142 nsew signal output
rlabel metal2 s 51814 193832 51870 194632 6 d_out[32]
port 143 nsew signal output
rlabel metal2 s 52734 193832 52790 194632 6 d_out[33]
port 144 nsew signal output
rlabel metal2 s 53654 193832 53710 194632 6 d_out[34]
port 145 nsew signal output
rlabel metal2 s 54482 193832 54538 194632 6 d_out[35]
port 146 nsew signal output
rlabel metal2 s 55402 193832 55458 194632 6 d_out[36]
port 147 nsew signal output
rlabel metal2 s 56322 193832 56378 194632 6 d_out[37]
port 148 nsew signal output
rlabel metal2 s 57242 193832 57298 194632 6 d_out[38]
port 149 nsew signal output
rlabel metal2 s 58162 193832 58218 194632 6 d_out[39]
port 150 nsew signal output
rlabel metal2 s 25594 193832 25650 194632 6 d_out[3]
port 151 nsew signal output
rlabel metal2 s 59082 193832 59138 194632 6 d_out[40]
port 152 nsew signal output
rlabel metal2 s 59910 193832 59966 194632 6 d_out[41]
port 153 nsew signal output
rlabel metal2 s 60830 193832 60886 194632 6 d_out[42]
port 154 nsew signal output
rlabel metal2 s 61750 193832 61806 194632 6 d_out[43]
port 155 nsew signal output
rlabel metal2 s 62670 193832 62726 194632 6 d_out[44]
port 156 nsew signal output
rlabel metal2 s 63590 193832 63646 194632 6 d_out[45]
port 157 nsew signal output
rlabel metal2 s 64418 193832 64474 194632 6 d_out[46]
port 158 nsew signal output
rlabel metal2 s 65338 193832 65394 194632 6 d_out[47]
port 159 nsew signal output
rlabel metal2 s 66258 193832 66314 194632 6 d_out[48]
port 160 nsew signal output
rlabel metal2 s 67178 193832 67234 194632 6 d_out[49]
port 161 nsew signal output
rlabel metal2 s 26514 193832 26570 194632 6 d_out[4]
port 162 nsew signal output
rlabel metal2 s 68098 193832 68154 194632 6 d_out[50]
port 163 nsew signal output
rlabel metal2 s 68926 193832 68982 194632 6 d_out[51]
port 164 nsew signal output
rlabel metal2 s 69846 193832 69902 194632 6 d_out[52]
port 165 nsew signal output
rlabel metal2 s 70766 193832 70822 194632 6 d_out[53]
port 166 nsew signal output
rlabel metal2 s 71686 193832 71742 194632 6 d_out[54]
port 167 nsew signal output
rlabel metal2 s 72606 193832 72662 194632 6 d_out[55]
port 168 nsew signal output
rlabel metal2 s 73526 193832 73582 194632 6 d_out[56]
port 169 nsew signal output
rlabel metal2 s 74354 193832 74410 194632 6 d_out[57]
port 170 nsew signal output
rlabel metal2 s 75274 193832 75330 194632 6 d_out[58]
port 171 nsew signal output
rlabel metal2 s 76194 193832 76250 194632 6 d_out[59]
port 172 nsew signal output
rlabel metal2 s 27434 193832 27490 194632 6 d_out[5]
port 173 nsew signal output
rlabel metal2 s 77114 193832 77170 194632 6 d_out[60]
port 174 nsew signal output
rlabel metal2 s 78034 193832 78090 194632 6 d_out[61]
port 175 nsew signal output
rlabel metal2 s 78862 193832 78918 194632 6 d_out[62]
port 176 nsew signal output
rlabel metal2 s 79782 193832 79838 194632 6 d_out[63]
port 177 nsew signal output
rlabel metal2 s 80702 193832 80758 194632 6 d_out[64]
port 178 nsew signal output
rlabel metal2 s 81622 193832 81678 194632 6 d_out[65]
port 179 nsew signal output
rlabel metal2 s 82542 193832 82598 194632 6 d_out[66]
port 180 nsew signal output
rlabel metal2 s 83462 193832 83518 194632 6 d_out[67]
port 181 nsew signal output
rlabel metal2 s 84290 193832 84346 194632 6 d_out[68]
port 182 nsew signal output
rlabel metal2 s 85210 193832 85266 194632 6 d_out[69]
port 183 nsew signal output
rlabel metal2 s 28354 193832 28410 194632 6 d_out[6]
port 184 nsew signal output
rlabel metal2 s 86130 193832 86186 194632 6 d_out[70]
port 185 nsew signal output
rlabel metal2 s 87050 193832 87106 194632 6 d_out[71]
port 186 nsew signal output
rlabel metal2 s 87970 193832 88026 194632 6 d_out[72]
port 187 nsew signal output
rlabel metal2 s 88798 193832 88854 194632 6 d_out[73]
port 188 nsew signal output
rlabel metal2 s 89718 193832 89774 194632 6 d_out[74]
port 189 nsew signal output
rlabel metal2 s 90638 193832 90694 194632 6 d_out[75]
port 190 nsew signal output
rlabel metal2 s 91558 193832 91614 194632 6 d_out[76]
port 191 nsew signal output
rlabel metal2 s 92478 193832 92534 194632 6 d_out[77]
port 192 nsew signal output
rlabel metal2 s 93398 193832 93454 194632 6 d_out[78]
port 193 nsew signal output
rlabel metal2 s 94226 193832 94282 194632 6 d_out[79]
port 194 nsew signal output
rlabel metal2 s 29274 193832 29330 194632 6 d_out[7]
port 195 nsew signal output
rlabel metal2 s 95146 193832 95202 194632 6 d_out[80]
port 196 nsew signal output
rlabel metal2 s 96066 193832 96122 194632 6 d_out[81]
port 197 nsew signal output
rlabel metal2 s 96986 193832 97042 194632 6 d_out[82]
port 198 nsew signal output
rlabel metal2 s 97906 193832 97962 194632 6 d_out[83]
port 199 nsew signal output
rlabel metal2 s 98734 193832 98790 194632 6 d_out[84]
port 200 nsew signal output
rlabel metal2 s 99654 193832 99710 194632 6 d_out[85]
port 201 nsew signal output
rlabel metal2 s 100574 193832 100630 194632 6 d_out[86]
port 202 nsew signal output
rlabel metal2 s 101494 193832 101550 194632 6 d_out[87]
port 203 nsew signal output
rlabel metal2 s 102414 193832 102470 194632 6 d_out[88]
port 204 nsew signal output
rlabel metal2 s 103242 193832 103298 194632 6 d_out[89]
port 205 nsew signal output
rlabel metal2 s 30102 193832 30158 194632 6 d_out[8]
port 206 nsew signal output
rlabel metal2 s 104162 193832 104218 194632 6 d_out[90]
port 207 nsew signal output
rlabel metal2 s 105082 193832 105138 194632 6 d_out[91]
port 208 nsew signal output
rlabel metal2 s 106002 193832 106058 194632 6 d_out[92]
port 209 nsew signal output
rlabel metal2 s 106922 193832 106978 194632 6 d_out[93]
port 210 nsew signal output
rlabel metal2 s 107842 193832 107898 194632 6 d_out[94]
port 211 nsew signal output
rlabel metal2 s 108670 193832 108726 194632 6 d_out[95]
port 212 nsew signal output
rlabel metal2 s 109590 193832 109646 194632 6 d_out[96]
port 213 nsew signal output
rlabel metal2 s 110510 193832 110566 194632 6 d_out[97]
port 214 nsew signal output
rlabel metal2 s 111430 193832 111486 194632 6 d_out[98]
port 215 nsew signal output
rlabel metal2 s 112350 193832 112406 194632 6 d_out[99]
port 216 nsew signal output
rlabel metal2 s 31022 193832 31078 194632 6 d_out[9]
port 217 nsew signal output
rlabel metal3 s 0 0 800 120 6 w_in[0]
port 218 nsew signal input
rlabel metal3 s 0 27200 800 27320 6 w_in[10]
port 219 nsew signal input
rlabel metal3 s 0 29920 800 30040 6 w_in[11]
port 220 nsew signal input
rlabel metal3 s 0 32640 800 32760 6 w_in[12]
port 221 nsew signal input
rlabel metal3 s 0 35360 800 35480 6 w_in[13]
port 222 nsew signal input
rlabel metal3 s 0 38080 800 38200 6 w_in[14]
port 223 nsew signal input
rlabel metal3 s 0 40800 800 40920 6 w_in[15]
port 224 nsew signal input
rlabel metal3 s 0 43520 800 43640 6 w_in[16]
port 225 nsew signal input
rlabel metal3 s 0 46240 800 46360 6 w_in[17]
port 226 nsew signal input
rlabel metal3 s 0 48960 800 49080 6 w_in[18]
port 227 nsew signal input
rlabel metal3 s 0 51680 800 51800 6 w_in[19]
port 228 nsew signal input
rlabel metal3 s 0 2720 800 2840 6 w_in[1]
port 229 nsew signal input
rlabel metal3 s 0 54400 800 54520 6 w_in[20]
port 230 nsew signal input
rlabel metal3 s 0 57120 800 57240 6 w_in[21]
port 231 nsew signal input
rlabel metal3 s 0 59840 800 59960 6 w_in[22]
port 232 nsew signal input
rlabel metal3 s 0 62560 800 62680 6 w_in[23]
port 233 nsew signal input
rlabel metal3 s 0 65280 800 65400 6 w_in[24]
port 234 nsew signal input
rlabel metal3 s 0 68000 800 68120 6 w_in[25]
port 235 nsew signal input
rlabel metal3 s 0 70720 800 70840 6 w_in[26]
port 236 nsew signal input
rlabel metal3 s 0 73440 800 73560 6 w_in[27]
port 237 nsew signal input
rlabel metal3 s 0 76160 800 76280 6 w_in[28]
port 238 nsew signal input
rlabel metal3 s 0 78880 800 79000 6 w_in[29]
port 239 nsew signal input
rlabel metal3 s 0 5440 800 5560 6 w_in[2]
port 240 nsew signal input
rlabel metal3 s 0 81600 800 81720 6 w_in[30]
port 241 nsew signal input
rlabel metal3 s 0 84320 800 84440 6 w_in[31]
port 242 nsew signal input
rlabel metal3 s 0 87040 800 87160 6 w_in[32]
port 243 nsew signal input
rlabel metal3 s 0 89760 800 89880 6 w_in[33]
port 244 nsew signal input
rlabel metal3 s 0 92480 800 92600 6 w_in[34]
port 245 nsew signal input
rlabel metal3 s 0 95200 800 95320 6 w_in[35]
port 246 nsew signal input
rlabel metal3 s 0 97920 800 98040 6 w_in[36]
port 247 nsew signal input
rlabel metal3 s 0 100640 800 100760 6 w_in[37]
port 248 nsew signal input
rlabel metal3 s 0 103360 800 103480 6 w_in[38]
port 249 nsew signal input
rlabel metal3 s 0 106080 800 106200 6 w_in[39]
port 250 nsew signal input
rlabel metal3 s 0 8160 800 8280 6 w_in[3]
port 251 nsew signal input
rlabel metal3 s 0 108800 800 108920 6 w_in[40]
port 252 nsew signal input
rlabel metal3 s 0 111520 800 111640 6 w_in[41]
port 253 nsew signal input
rlabel metal3 s 0 114240 800 114360 6 w_in[42]
port 254 nsew signal input
rlabel metal3 s 0 116960 800 117080 6 w_in[43]
port 255 nsew signal input
rlabel metal3 s 0 119680 800 119800 6 w_in[44]
port 256 nsew signal input
rlabel metal3 s 0 122400 800 122520 6 w_in[45]
port 257 nsew signal input
rlabel metal3 s 0 125120 800 125240 6 w_in[46]
port 258 nsew signal input
rlabel metal3 s 0 127840 800 127960 6 w_in[47]
port 259 nsew signal input
rlabel metal3 s 0 130560 800 130680 6 w_in[48]
port 260 nsew signal input
rlabel metal3 s 0 133280 800 133400 6 w_in[49]
port 261 nsew signal input
rlabel metal3 s 0 10880 800 11000 6 w_in[4]
port 262 nsew signal input
rlabel metal3 s 0 136000 800 136120 6 w_in[50]
port 263 nsew signal input
rlabel metal3 s 0 138720 800 138840 6 w_in[51]
port 264 nsew signal input
rlabel metal3 s 0 141440 800 141560 6 w_in[52]
port 265 nsew signal input
rlabel metal3 s 0 144160 800 144280 6 w_in[53]
port 266 nsew signal input
rlabel metal3 s 0 146880 800 147000 6 w_in[54]
port 267 nsew signal input
rlabel metal3 s 0 149600 800 149720 6 w_in[55]
port 268 nsew signal input
rlabel metal3 s 0 152320 800 152440 6 w_in[56]
port 269 nsew signal input
rlabel metal3 s 0 155040 800 155160 6 w_in[57]
port 270 nsew signal input
rlabel metal3 s 0 157760 800 157880 6 w_in[58]
port 271 nsew signal input
rlabel metal3 s 0 160480 800 160600 6 w_in[59]
port 272 nsew signal input
rlabel metal3 s 0 13600 800 13720 6 w_in[5]
port 273 nsew signal input
rlabel metal3 s 0 163200 800 163320 6 w_in[60]
port 274 nsew signal input
rlabel metal3 s 0 165920 800 166040 6 w_in[61]
port 275 nsew signal input
rlabel metal3 s 0 168640 800 168760 6 w_in[62]
port 276 nsew signal input
rlabel metal3 s 0 171360 800 171480 6 w_in[63]
port 277 nsew signal input
rlabel metal3 s 0 174080 800 174200 6 w_in[64]
port 278 nsew signal input
rlabel metal3 s 0 176800 800 176920 6 w_in[65]
port 279 nsew signal input
rlabel metal3 s 0 179520 800 179640 6 w_in[66]
port 280 nsew signal input
rlabel metal3 s 0 182240 800 182360 6 w_in[67]
port 281 nsew signal input
rlabel metal3 s 0 184960 800 185080 6 w_in[68]
port 282 nsew signal input
rlabel metal3 s 0 187680 800 187800 6 w_in[69]
port 283 nsew signal input
rlabel metal3 s 0 16320 800 16440 6 w_in[6]
port 284 nsew signal input
rlabel metal3 s 0 190400 800 190520 6 w_in[70]
port 285 nsew signal input
rlabel metal3 s 0 193120 800 193240 6 w_in[71]
port 286 nsew signal input
rlabel metal3 s 0 19040 800 19160 6 w_in[7]
port 287 nsew signal input
rlabel metal3 s 0 21760 800 21880 6 w_in[8]
port 288 nsew signal input
rlabel metal3 s 0 24480 800 24600 6 w_in[9]
port 289 nsew signal input
rlabel metal4 s 188528 760 188848 192344 6 vccd1
port 290 nsew power bidirectional
rlabel metal4 s 157808 760 158128 192344 6 vccd1
port 291 nsew power bidirectional
rlabel metal4 s 127088 760 127408 192344 6 vccd1
port 292 nsew power bidirectional
rlabel metal4 s 96368 760 96688 192344 6 vccd1
port 293 nsew power bidirectional
rlabel metal4 s 65648 760 65968 192344 6 vccd1
port 294 nsew power bidirectional
rlabel metal4 s 34928 760 35248 192344 6 vccd1
port 295 nsew power bidirectional
rlabel metal4 s 4208 760 4528 192344 6 vccd1
port 296 nsew power bidirectional
rlabel metal4 s 173168 760 173488 192344 6 vssd1
port 297 nsew ground bidirectional
rlabel metal4 s 142448 760 142768 192344 6 vssd1
port 298 nsew ground bidirectional
rlabel metal4 s 111728 760 112048 192344 6 vssd1
port 299 nsew ground bidirectional
rlabel metal4 s 81008 760 81328 192344 6 vssd1
port 300 nsew ground bidirectional
rlabel metal4 s 50288 760 50608 192344 6 vssd1
port 301 nsew ground bidirectional
rlabel metal4 s 19568 760 19888 192344 6 vssd1
port 302 nsew ground bidirectional
rlabel metal4 s 189188 808 189508 192296 6 vccd2
port 303 nsew power bidirectional
rlabel metal4 s 158468 808 158788 192296 6 vccd2
port 304 nsew power bidirectional
rlabel metal4 s 127748 808 128068 192296 6 vccd2
port 305 nsew power bidirectional
rlabel metal4 s 97028 808 97348 192296 6 vccd2
port 306 nsew power bidirectional
rlabel metal4 s 66308 808 66628 192296 6 vccd2
port 307 nsew power bidirectional
rlabel metal4 s 35588 808 35908 192296 6 vccd2
port 308 nsew power bidirectional
rlabel metal4 s 4868 808 5188 192296 6 vccd2
port 309 nsew power bidirectional
rlabel metal4 s 173828 808 174148 192296 6 vssd2
port 310 nsew ground bidirectional
rlabel metal4 s 143108 808 143428 192296 6 vssd2
port 311 nsew ground bidirectional
rlabel metal4 s 112388 808 112708 192296 6 vssd2
port 312 nsew ground bidirectional
rlabel metal4 s 81668 808 81988 192296 6 vssd2
port 313 nsew ground bidirectional
rlabel metal4 s 50948 808 51268 192296 6 vssd2
port 314 nsew ground bidirectional
rlabel metal4 s 20228 808 20548 192296 6 vssd2
port 315 nsew ground bidirectional
rlabel metal4 s 189848 808 190168 192296 6 vdda1
port 316 nsew power bidirectional
rlabel metal4 s 159128 808 159448 192296 6 vdda1
port 317 nsew power bidirectional
rlabel metal4 s 128408 808 128728 192296 6 vdda1
port 318 nsew power bidirectional
rlabel metal4 s 97688 808 98008 192296 6 vdda1
port 319 nsew power bidirectional
rlabel metal4 s 66968 808 67288 192296 6 vdda1
port 320 nsew power bidirectional
rlabel metal4 s 36248 808 36568 192296 6 vdda1
port 321 nsew power bidirectional
rlabel metal4 s 5528 808 5848 192296 6 vdda1
port 322 nsew power bidirectional
rlabel metal4 s 174488 808 174808 192296 6 vssa1
port 323 nsew ground bidirectional
rlabel metal4 s 143768 808 144088 192296 6 vssa1
port 324 nsew ground bidirectional
rlabel metal4 s 113048 808 113368 192296 6 vssa1
port 325 nsew ground bidirectional
rlabel metal4 s 82328 808 82648 192296 6 vssa1
port 326 nsew ground bidirectional
rlabel metal4 s 51608 808 51928 192296 6 vssa1
port 327 nsew ground bidirectional
rlabel metal4 s 20888 808 21208 192296 6 vssa1
port 328 nsew ground bidirectional
rlabel metal4 s 190508 808 190828 192296 6 vdda2
port 329 nsew power bidirectional
rlabel metal4 s 159788 808 160108 192296 6 vdda2
port 330 nsew power bidirectional
rlabel metal4 s 129068 808 129388 192296 6 vdda2
port 331 nsew power bidirectional
rlabel metal4 s 98348 808 98668 192296 6 vdda2
port 332 nsew power bidirectional
rlabel metal4 s 67628 808 67948 192296 6 vdda2
port 333 nsew power bidirectional
rlabel metal4 s 36908 808 37228 192296 6 vdda2
port 334 nsew power bidirectional
rlabel metal4 s 6188 808 6508 192296 6 vdda2
port 335 nsew power bidirectional
rlabel metal4 s 175148 808 175468 192296 6 vssa2
port 336 nsew ground bidirectional
rlabel metal4 s 144428 808 144748 192296 6 vssa2
port 337 nsew ground bidirectional
rlabel metal4 s 113708 808 114028 192296 6 vssa2
port 338 nsew ground bidirectional
rlabel metal4 s 82988 808 83308 192296 6 vssa2
port 339 nsew ground bidirectional
rlabel metal4 s 52268 808 52588 192296 6 vssa2
port 340 nsew ground bidirectional
rlabel metal4 s 21548 808 21868 192296 6 vssa2
port 341 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 195482 194632
string LEFview TRUE
<< end >>
