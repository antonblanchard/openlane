VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM_512x64
  CLASS BLOCK ;
  FOREIGN RAM_512x64 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2788.900 BY 789.040 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2441.960 0.000 2442.240 4.000 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2460.820 0.000 2461.100 4.000 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2480.140 0.000 2480.420 4.000 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2499.000 0.000 2499.280 4.000 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2517.860 0.000 2518.140 4.000 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2537.180 0.000 2537.460 4.000 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2556.040 0.000 2556.320 4.000 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2575.360 0.000 2575.640 4.000 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2594.220 0.000 2594.500 4.000 ;
    END
  END A[8]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2613.080 0.000 2613.360 4.000 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1222.960 0.000 1223.240 4.000 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.400 0.000 1413.680 4.000 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.260 0.000 1432.540 4.000 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1451.580 0.000 1451.860 4.000 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1470.440 0.000 1470.720 4.000 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.300 0.000 1489.580 4.000 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1508.620 0.000 1508.900 4.000 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.480 0.000 1527.760 4.000 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1546.800 0.000 1547.080 4.000 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.660 0.000 1565.940 4.000 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.520 0.000 1584.800 4.000 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1241.820 0.000 1242.100 4.000 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.840 0.000 1604.120 4.000 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.700 0.000 1622.980 4.000 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1642.020 0.000 1642.300 4.000 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1660.880 0.000 1661.160 4.000 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.740 0.000 1680.020 4.000 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.060 0.000 1699.340 4.000 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1717.920 0.000 1718.200 4.000 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1737.240 0.000 1737.520 4.000 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1756.100 0.000 1756.380 4.000 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.960 0.000 1775.240 4.000 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.680 0.000 1260.960 4.000 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1794.280 0.000 1794.560 4.000 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1813.140 0.000 1813.420 4.000 ;
    END
  END Di[31]
  PIN Di[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1832.460 0.000 1832.740 4.000 ;
    END
  END Di[32]
  PIN Di[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1851.320 0.000 1851.600 4.000 ;
    END
  END Di[33]
  PIN Di[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.640 0.000 1870.920 4.000 ;
    END
  END Di[34]
  PIN Di[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1889.500 0.000 1889.780 4.000 ;
    END
  END Di[35]
  PIN Di[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1908.360 0.000 1908.640 4.000 ;
    END
  END Di[36]
  PIN Di[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1927.680 0.000 1927.960 4.000 ;
    END
  END Di[37]
  PIN Di[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1946.540 0.000 1946.820 4.000 ;
    END
  END Di[38]
  PIN Di[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.860 0.000 1966.140 4.000 ;
    END
  END Di[39]
  PIN Di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.000 0.000 1280.280 4.000 ;
    END
  END Di[3]
  PIN Di[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1984.720 0.000 1985.000 4.000 ;
    END
  END Di[40]
  PIN Di[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2003.580 0.000 2003.860 4.000 ;
    END
  END Di[41]
  PIN Di[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2022.900 0.000 2023.180 4.000 ;
    END
  END Di[42]
  PIN Di[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.760 0.000 2042.040 4.000 ;
    END
  END Di[43]
  PIN Di[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2061.080 0.000 2061.360 4.000 ;
    END
  END Di[44]
  PIN Di[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2079.940 0.000 2080.220 4.000 ;
    END
  END Di[45]
  PIN Di[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2098.800 0.000 2099.080 4.000 ;
    END
  END Di[46]
  PIN Di[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.120 0.000 2118.400 4.000 ;
    END
  END Di[47]
  PIN Di[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.980 0.000 2137.260 4.000 ;
    END
  END Di[48]
  PIN Di[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2156.300 0.000 2156.580 4.000 ;
    END
  END Di[49]
  PIN Di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.860 0.000 1299.140 4.000 ;
    END
  END Di[4]
  PIN Di[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2175.160 0.000 2175.440 4.000 ;
    END
  END Di[50]
  PIN Di[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2194.020 0.000 2194.300 4.000 ;
    END
  END Di[51]
  PIN Di[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.340 0.000 2213.620 4.000 ;
    END
  END Di[52]
  PIN Di[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2232.200 0.000 2232.480 4.000 ;
    END
  END Di[53]
  PIN Di[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2251.520 0.000 2251.800 4.000 ;
    END
  END Di[54]
  PIN Di[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2270.380 0.000 2270.660 4.000 ;
    END
  END Di[55]
  PIN Di[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2289.240 0.000 2289.520 4.000 ;
    END
  END Di[56]
  PIN Di[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2308.560 0.000 2308.840 4.000 ;
    END
  END Di[57]
  PIN Di[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2327.420 0.000 2327.700 4.000 ;
    END
  END Di[58]
  PIN Di[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2346.740 0.000 2347.020 4.000 ;
    END
  END Di[59]
  PIN Di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1318.180 0.000 1318.460 4.000 ;
    END
  END Di[5]
  PIN Di[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2365.600 0.000 2365.880 4.000 ;
    END
  END Di[60]
  PIN Di[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.920 0.000 2385.200 4.000 ;
    END
  END Di[61]
  PIN Di[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2403.780 0.000 2404.060 4.000 ;
    END
  END Di[62]
  PIN Di[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2422.640 0.000 2422.920 4.000 ;
    END
  END Di[63]
  PIN Di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1337.040 0.000 1337.320 4.000 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.900 0.000 1356.180 4.000 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.220 0.000 1375.500 4.000 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.080 0.000 1394.360 4.000 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.960 0.000 4.240 4.000 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.400 0.000 194.680 4.000 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.260 0.000 213.540 4.000 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.120 0.000 232.400 4.000 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.440 0.000 251.720 4.000 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.300 0.000 270.580 4.000 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.620 0.000 289.900 4.000 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.480 0.000 308.760 4.000 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.340 0.000 327.620 4.000 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.660 0.000 346.940 4.000 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.520 0.000 365.800 4.000 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.820 0.000 23.100 4.000 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.840 0.000 385.120 4.000 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.700 0.000 403.980 4.000 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.560 0.000 422.840 4.000 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.880 0.000 442.160 4.000 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.740 0.000 461.020 4.000 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.060 0.000 480.340 4.000 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.920 0.000 499.200 4.000 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.240 0.000 518.520 4.000 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.100 0.000 537.380 4.000 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.960 0.000 556.240 4.000 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.680 0.000 41.960 4.000 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.280 0.000 575.560 4.000 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.140 0.000 594.420 4.000 ;
    END
  END Do[31]
  PIN Do[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.460 0.000 613.740 4.000 ;
    END
  END Do[32]
  PIN Do[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.320 0.000 632.600 4.000 ;
    END
  END Do[33]
  PIN Do[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.180 0.000 651.460 4.000 ;
    END
  END Do[34]
  PIN Do[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.500 0.000 670.780 4.000 ;
    END
  END Do[35]
  PIN Do[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.360 0.000 689.640 4.000 ;
    END
  END Do[36]
  PIN Do[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.680 0.000 708.960 4.000 ;
    END
  END Do[37]
  PIN Do[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.540 0.000 727.820 4.000 ;
    END
  END Do[38]
  PIN Do[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.400 0.000 746.680 4.000 ;
    END
  END Do[39]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.000 0.000 61.280 4.000 ;
    END
  END Do[3]
  PIN Do[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.720 0.000 766.000 4.000 ;
    END
  END Do[40]
  PIN Do[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.580 0.000 784.860 4.000 ;
    END
  END Do[41]
  PIN Do[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.900 0.000 804.180 4.000 ;
    END
  END Do[42]
  PIN Do[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.760 0.000 823.040 4.000 ;
    END
  END Do[43]
  PIN Do[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.620 0.000 841.900 4.000 ;
    END
  END Do[44]
  PIN Do[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.940 0.000 861.220 4.000 ;
    END
  END Do[45]
  PIN Do[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.800 0.000 880.080 4.000 ;
    END
  END Do[46]
  PIN Do[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.120 0.000 899.400 4.000 ;
    END
  END Do[47]
  PIN Do[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.980 0.000 918.260 4.000 ;
    END
  END Do[48]
  PIN Do[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.300 0.000 937.580 4.000 ;
    END
  END Do[49]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.860 0.000 80.140 4.000 ;
    END
  END Do[4]
  PIN Do[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.160 0.000 956.440 4.000 ;
    END
  END Do[50]
  PIN Do[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.020 0.000 975.300 4.000 ;
    END
  END Do[51]
  PIN Do[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.340 0.000 994.620 4.000 ;
    END
  END Do[52]
  PIN Do[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.200 0.000 1013.480 4.000 ;
    END
  END Do[53]
  PIN Do[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1032.520 0.000 1032.800 4.000 ;
    END
  END Do[54]
  PIN Do[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.380 0.000 1051.660 4.000 ;
    END
  END Do[55]
  PIN Do[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.240 0.000 1070.520 4.000 ;
    END
  END Do[56]
  PIN Do[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1089.560 0.000 1089.840 4.000 ;
    END
  END Do[57]
  PIN Do[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.420 0.000 1108.700 4.000 ;
    END
  END Do[58]
  PIN Do[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.740 0.000 1128.020 4.000 ;
    END
  END Do[59]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.180 0.000 99.460 4.000 ;
    END
  END Do[5]
  PIN Do[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.600 0.000 1146.880 4.000 ;
    END
  END Do[60]
  PIN Do[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.460 0.000 1165.740 4.000 ;
    END
  END Do[61]
  PIN Do[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.780 0.000 1185.060 4.000 ;
    END
  END Do[62]
  PIN Do[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.640 0.000 1203.920 4.000 ;
    END
  END Do[63]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.040 0.000 118.320 4.000 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.900 0.000 137.180 4.000 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.220 0.000 156.500 4.000 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.080 0.000 175.360 4.000 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2784.660 0.000 2784.940 4.000 ;
    END
  END EN
  PIN WE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.400 0.000 2632.680 4.000 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2651.260 0.000 2651.540 4.000 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2670.580 0.000 2670.860 4.000 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2689.440 0.000 2689.720 4.000 ;
    END
  END WE[3]
  PIN WE[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2708.300 0.000 2708.580 4.000 ;
    END
  END WE[4]
  PIN WE[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2727.620 0.000 2727.900 4.000 ;
    END
  END WE[5]
  PIN WE[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2746.480 0.000 2746.760 4.000 ;
    END
  END WE[6]
  PIN WE[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2765.800 0.000 2766.080 4.000 ;
    END
  END WE[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2780.510 10.640 2782.110 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2626.910 10.640 2628.510 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2473.310 10.640 2474.910 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2319.710 10.640 2321.310 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2166.110 10.640 2167.710 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2012.510 10.640 2014.110 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1858.910 10.640 1860.510 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1705.310 10.640 1706.910 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1551.710 10.640 1553.310 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1398.110 10.640 1399.710 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1244.510 10.640 1246.110 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1090.910 10.640 1092.510 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 937.310 10.640 938.910 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 783.710 10.640 785.310 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 630.110 10.640 631.710 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 476.510 10.640 478.110 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 322.910 10.640 324.510 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 169.310 10.640 170.910 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.710 10.640 17.310 789.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2703.710 10.640 2705.310 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2550.110 10.640 2551.710 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2396.510 10.640 2398.110 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2242.910 10.640 2244.510 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2089.310 10.640 2090.910 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1935.710 10.640 1937.310 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1782.110 10.640 1783.710 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1628.510 10.640 1630.110 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1474.910 10.640 1476.510 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1321.310 10.640 1322.910 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1167.710 10.640 1169.310 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1014.110 10.640 1015.710 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 860.510 10.640 862.110 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 706.910 10.640 708.510 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 553.310 10.640 554.910 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 399.710 10.640 401.310 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 246.110 10.640 247.710 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 92.510 10.640 94.110 789.040 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2783.810 10.880 2785.410 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2630.210 10.880 2631.810 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2476.610 10.880 2478.210 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2323.010 10.880 2324.610 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2169.410 10.880 2171.010 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2015.810 10.880 2017.410 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1862.210 10.880 1863.810 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1708.610 10.880 1710.210 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1555.010 10.880 1556.610 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1401.410 10.880 1403.010 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1247.810 10.880 1249.410 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1094.210 10.880 1095.810 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 940.610 10.880 942.210 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 787.010 10.880 788.610 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 633.410 10.880 635.010 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 479.810 10.880 481.410 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 326.210 10.880 327.810 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 172.610 10.880 174.210 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.010 10.880 20.610 788.800 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2707.010 10.880 2708.610 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2553.410 10.880 2555.010 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2399.810 10.880 2401.410 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2246.210 10.880 2247.810 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2092.610 10.880 2094.210 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1939.010 10.880 1940.610 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1785.410 10.880 1787.010 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1631.810 10.880 1633.410 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1478.210 10.880 1479.810 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1324.610 10.880 1326.210 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1171.010 10.880 1172.610 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1017.410 10.880 1019.010 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 863.810 10.880 865.410 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 710.210 10.880 711.810 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 556.610 10.880 558.210 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 403.010 10.880 404.610 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 249.410 10.880 251.010 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.810 10.880 97.410 788.800 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2633.510 10.880 2635.110 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2479.910 10.880 2481.510 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2326.310 10.880 2327.910 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2172.710 10.880 2174.310 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2019.110 10.880 2020.710 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1865.510 10.880 1867.110 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1711.910 10.880 1713.510 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1558.310 10.880 1559.910 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1404.710 10.880 1406.310 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1251.110 10.880 1252.710 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1097.510 10.880 1099.110 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 943.910 10.880 945.510 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 790.310 10.880 791.910 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 636.710 10.880 638.310 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 483.110 10.880 484.710 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 329.510 10.880 331.110 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 175.910 10.880 177.510 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.310 10.880 23.910 788.800 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2710.310 10.880 2711.910 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2556.710 10.880 2558.310 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2403.110 10.880 2404.710 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2249.510 10.880 2251.110 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2095.910 10.880 2097.510 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1942.310 10.880 1943.910 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1788.710 10.880 1790.310 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1635.110 10.880 1636.710 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1481.510 10.880 1483.110 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1327.910 10.880 1329.510 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1174.310 10.880 1175.910 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1020.710 10.880 1022.310 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 867.110 10.880 868.710 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 713.510 10.880 715.110 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 559.910 10.880 561.510 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 406.310 10.880 407.910 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 252.710 10.880 254.310 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 99.110 10.880 100.710 788.800 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2636.810 10.880 2638.410 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2483.210 10.880 2484.810 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2329.610 10.880 2331.210 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2176.010 10.880 2177.610 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2022.410 10.880 2024.010 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1868.810 10.880 1870.410 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1715.210 10.880 1716.810 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1561.610 10.880 1563.210 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1408.010 10.880 1409.610 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1254.410 10.880 1256.010 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1100.810 10.880 1102.410 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 947.210 10.880 948.810 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 793.610 10.880 795.210 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 640.010 10.880 641.610 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 486.410 10.880 488.010 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 332.810 10.880 334.410 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 179.210 10.880 180.810 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 25.610 10.880 27.210 788.800 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2713.610 10.880 2715.210 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2560.010 10.880 2561.610 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2406.410 10.880 2408.010 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2252.810 10.880 2254.410 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2099.210 10.880 2100.810 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1945.610 10.880 1947.210 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1792.010 10.880 1793.610 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1638.410 10.880 1640.010 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1484.810 10.880 1486.410 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1331.210 10.880 1332.810 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1177.610 10.880 1179.210 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1024.010 10.880 1025.610 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 870.410 10.880 872.010 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 716.810 10.880 718.410 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 563.210 10.880 564.810 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 409.610 10.880 411.210 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 256.010 10.880 257.610 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 102.410 10.880 104.010 788.800 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 0.190 6.545 2788.710 788.885 ;
      LAYER met1 ;
        RECT 0.190 6.500 2788.710 789.040 ;
      LAYER met2 ;
        RECT 2.590 4.280 2786.770 789.040 ;
        RECT 2.590 4.000 3.680 4.280 ;
        RECT 4.520 4.000 22.540 4.280 ;
        RECT 23.380 4.000 41.400 4.280 ;
        RECT 42.240 4.000 60.720 4.280 ;
        RECT 61.560 4.000 79.580 4.280 ;
        RECT 80.420 4.000 98.900 4.280 ;
        RECT 99.740 4.000 117.760 4.280 ;
        RECT 118.600 4.000 136.620 4.280 ;
        RECT 137.460 4.000 155.940 4.280 ;
        RECT 156.780 4.000 174.800 4.280 ;
        RECT 175.640 4.000 194.120 4.280 ;
        RECT 194.960 4.000 212.980 4.280 ;
        RECT 213.820 4.000 231.840 4.280 ;
        RECT 232.680 4.000 251.160 4.280 ;
        RECT 252.000 4.000 270.020 4.280 ;
        RECT 270.860 4.000 289.340 4.280 ;
        RECT 290.180 4.000 308.200 4.280 ;
        RECT 309.040 4.000 327.060 4.280 ;
        RECT 327.900 4.000 346.380 4.280 ;
        RECT 347.220 4.000 365.240 4.280 ;
        RECT 366.080 4.000 384.560 4.280 ;
        RECT 385.400 4.000 403.420 4.280 ;
        RECT 404.260 4.000 422.280 4.280 ;
        RECT 423.120 4.000 441.600 4.280 ;
        RECT 442.440 4.000 460.460 4.280 ;
        RECT 461.300 4.000 479.780 4.280 ;
        RECT 480.620 4.000 498.640 4.280 ;
        RECT 499.480 4.000 517.960 4.280 ;
        RECT 518.800 4.000 536.820 4.280 ;
        RECT 537.660 4.000 555.680 4.280 ;
        RECT 556.520 4.000 575.000 4.280 ;
        RECT 575.840 4.000 593.860 4.280 ;
        RECT 594.700 4.000 613.180 4.280 ;
        RECT 614.020 4.000 632.040 4.280 ;
        RECT 632.880 4.000 650.900 4.280 ;
        RECT 651.740 4.000 670.220 4.280 ;
        RECT 671.060 4.000 689.080 4.280 ;
        RECT 689.920 4.000 708.400 4.280 ;
        RECT 709.240 4.000 727.260 4.280 ;
        RECT 728.100 4.000 746.120 4.280 ;
        RECT 746.960 4.000 765.440 4.280 ;
        RECT 766.280 4.000 784.300 4.280 ;
        RECT 785.140 4.000 803.620 4.280 ;
        RECT 804.460 4.000 822.480 4.280 ;
        RECT 823.320 4.000 841.340 4.280 ;
        RECT 842.180 4.000 860.660 4.280 ;
        RECT 861.500 4.000 879.520 4.280 ;
        RECT 880.360 4.000 898.840 4.280 ;
        RECT 899.680 4.000 917.700 4.280 ;
        RECT 918.540 4.000 937.020 4.280 ;
        RECT 937.860 4.000 955.880 4.280 ;
        RECT 956.720 4.000 974.740 4.280 ;
        RECT 975.580 4.000 994.060 4.280 ;
        RECT 994.900 4.000 1012.920 4.280 ;
        RECT 1013.760 4.000 1032.240 4.280 ;
        RECT 1033.080 4.000 1051.100 4.280 ;
        RECT 1051.940 4.000 1069.960 4.280 ;
        RECT 1070.800 4.000 1089.280 4.280 ;
        RECT 1090.120 4.000 1108.140 4.280 ;
        RECT 1108.980 4.000 1127.460 4.280 ;
        RECT 1128.300 4.000 1146.320 4.280 ;
        RECT 1147.160 4.000 1165.180 4.280 ;
        RECT 1166.020 4.000 1184.500 4.280 ;
        RECT 1185.340 4.000 1203.360 4.280 ;
        RECT 1204.200 4.000 1222.680 4.280 ;
        RECT 1223.520 4.000 1241.540 4.280 ;
        RECT 1242.380 4.000 1260.400 4.280 ;
        RECT 1261.240 4.000 1279.720 4.280 ;
        RECT 1280.560 4.000 1298.580 4.280 ;
        RECT 1299.420 4.000 1317.900 4.280 ;
        RECT 1318.740 4.000 1336.760 4.280 ;
        RECT 1337.600 4.000 1355.620 4.280 ;
        RECT 1356.460 4.000 1374.940 4.280 ;
        RECT 1375.780 4.000 1393.800 4.280 ;
        RECT 1394.640 4.000 1413.120 4.280 ;
        RECT 1413.960 4.000 1431.980 4.280 ;
        RECT 1432.820 4.000 1451.300 4.280 ;
        RECT 1452.140 4.000 1470.160 4.280 ;
        RECT 1471.000 4.000 1489.020 4.280 ;
        RECT 1489.860 4.000 1508.340 4.280 ;
        RECT 1509.180 4.000 1527.200 4.280 ;
        RECT 1528.040 4.000 1546.520 4.280 ;
        RECT 1547.360 4.000 1565.380 4.280 ;
        RECT 1566.220 4.000 1584.240 4.280 ;
        RECT 1585.080 4.000 1603.560 4.280 ;
        RECT 1604.400 4.000 1622.420 4.280 ;
        RECT 1623.260 4.000 1641.740 4.280 ;
        RECT 1642.580 4.000 1660.600 4.280 ;
        RECT 1661.440 4.000 1679.460 4.280 ;
        RECT 1680.300 4.000 1698.780 4.280 ;
        RECT 1699.620 4.000 1717.640 4.280 ;
        RECT 1718.480 4.000 1736.960 4.280 ;
        RECT 1737.800 4.000 1755.820 4.280 ;
        RECT 1756.660 4.000 1774.680 4.280 ;
        RECT 1775.520 4.000 1794.000 4.280 ;
        RECT 1794.840 4.000 1812.860 4.280 ;
        RECT 1813.700 4.000 1832.180 4.280 ;
        RECT 1833.020 4.000 1851.040 4.280 ;
        RECT 1851.880 4.000 1870.360 4.280 ;
        RECT 1871.200 4.000 1889.220 4.280 ;
        RECT 1890.060 4.000 1908.080 4.280 ;
        RECT 1908.920 4.000 1927.400 4.280 ;
        RECT 1928.240 4.000 1946.260 4.280 ;
        RECT 1947.100 4.000 1965.580 4.280 ;
        RECT 1966.420 4.000 1984.440 4.280 ;
        RECT 1985.280 4.000 2003.300 4.280 ;
        RECT 2004.140 4.000 2022.620 4.280 ;
        RECT 2023.460 4.000 2041.480 4.280 ;
        RECT 2042.320 4.000 2060.800 4.280 ;
        RECT 2061.640 4.000 2079.660 4.280 ;
        RECT 2080.500 4.000 2098.520 4.280 ;
        RECT 2099.360 4.000 2117.840 4.280 ;
        RECT 2118.680 4.000 2136.700 4.280 ;
        RECT 2137.540 4.000 2156.020 4.280 ;
        RECT 2156.860 4.000 2174.880 4.280 ;
        RECT 2175.720 4.000 2193.740 4.280 ;
        RECT 2194.580 4.000 2213.060 4.280 ;
        RECT 2213.900 4.000 2231.920 4.280 ;
        RECT 2232.760 4.000 2251.240 4.280 ;
        RECT 2252.080 4.000 2270.100 4.280 ;
        RECT 2270.940 4.000 2288.960 4.280 ;
        RECT 2289.800 4.000 2308.280 4.280 ;
        RECT 2309.120 4.000 2327.140 4.280 ;
        RECT 2327.980 4.000 2346.460 4.280 ;
        RECT 2347.300 4.000 2365.320 4.280 ;
        RECT 2366.160 4.000 2384.640 4.280 ;
        RECT 2385.480 4.000 2403.500 4.280 ;
        RECT 2404.340 4.000 2422.360 4.280 ;
        RECT 2423.200 4.000 2441.680 4.280 ;
        RECT 2442.520 4.000 2460.540 4.280 ;
        RECT 2461.380 4.000 2479.860 4.280 ;
        RECT 2480.700 4.000 2498.720 4.280 ;
        RECT 2499.560 4.000 2517.580 4.280 ;
        RECT 2518.420 4.000 2536.900 4.280 ;
        RECT 2537.740 4.000 2555.760 4.280 ;
        RECT 2556.600 4.000 2575.080 4.280 ;
        RECT 2575.920 4.000 2593.940 4.280 ;
        RECT 2594.780 4.000 2612.800 4.280 ;
        RECT 2613.640 4.000 2632.120 4.280 ;
        RECT 2632.960 4.000 2650.980 4.280 ;
        RECT 2651.820 4.000 2670.300 4.280 ;
        RECT 2671.140 4.000 2689.160 4.280 ;
        RECT 2690.000 4.000 2708.020 4.280 ;
        RECT 2708.860 4.000 2727.340 4.280 ;
        RECT 2728.180 4.000 2746.200 4.280 ;
        RECT 2747.040 4.000 2765.520 4.280 ;
        RECT 2766.360 4.000 2784.380 4.280 ;
        RECT 2785.220 4.000 2786.770 4.280 ;
      LAYER met3 ;
        RECT 6.235 9.695 2785.885 788.965 ;
      LAYER met4 ;
        RECT 187.245 10.240 245.710 651.265 ;
        RECT 248.110 10.480 249.010 651.265 ;
        RECT 251.410 10.480 252.310 651.265 ;
        RECT 254.710 10.480 255.610 651.265 ;
        RECT 258.010 10.480 322.510 651.265 ;
        RECT 248.110 10.240 322.510 10.480 ;
        RECT 324.910 10.480 325.810 651.265 ;
        RECT 328.210 10.480 329.110 651.265 ;
        RECT 331.510 10.480 332.410 651.265 ;
        RECT 334.810 10.480 399.310 651.265 ;
        RECT 324.910 10.240 399.310 10.480 ;
        RECT 401.710 10.480 402.610 651.265 ;
        RECT 405.010 10.480 405.910 651.265 ;
        RECT 408.310 10.480 409.210 651.265 ;
        RECT 411.610 10.480 476.110 651.265 ;
        RECT 401.710 10.240 476.110 10.480 ;
        RECT 478.510 10.480 479.410 651.265 ;
        RECT 481.810 10.480 482.710 651.265 ;
        RECT 485.110 10.480 486.010 651.265 ;
        RECT 488.410 10.480 552.910 651.265 ;
        RECT 478.510 10.240 552.910 10.480 ;
        RECT 555.310 10.480 556.210 651.265 ;
        RECT 558.610 10.480 559.510 651.265 ;
        RECT 561.910 10.480 562.810 651.265 ;
        RECT 565.210 10.480 629.710 651.265 ;
        RECT 555.310 10.240 629.710 10.480 ;
        RECT 632.110 10.480 633.010 651.265 ;
        RECT 635.410 10.480 636.310 651.265 ;
        RECT 638.710 10.480 639.610 651.265 ;
        RECT 642.010 10.480 706.510 651.265 ;
        RECT 632.110 10.240 706.510 10.480 ;
        RECT 708.910 10.480 709.810 651.265 ;
        RECT 712.210 10.480 713.110 651.265 ;
        RECT 715.510 10.480 716.410 651.265 ;
        RECT 718.810 10.480 783.310 651.265 ;
        RECT 708.910 10.240 783.310 10.480 ;
        RECT 785.710 10.480 786.610 651.265 ;
        RECT 789.010 10.480 789.910 651.265 ;
        RECT 792.310 10.480 793.210 651.265 ;
        RECT 795.610 10.480 860.110 651.265 ;
        RECT 785.710 10.240 860.110 10.480 ;
        RECT 862.510 10.480 863.410 651.265 ;
        RECT 865.810 10.480 866.710 651.265 ;
        RECT 869.110 10.480 870.010 651.265 ;
        RECT 872.410 10.480 936.910 651.265 ;
        RECT 862.510 10.240 936.910 10.480 ;
        RECT 939.310 10.480 940.210 651.265 ;
        RECT 942.610 10.480 943.510 651.265 ;
        RECT 945.910 10.480 946.810 651.265 ;
        RECT 949.210 10.480 1013.710 651.265 ;
        RECT 939.310 10.240 1013.710 10.480 ;
        RECT 1016.110 10.480 1017.010 651.265 ;
        RECT 1019.410 10.480 1020.310 651.265 ;
        RECT 1022.710 10.480 1023.610 651.265 ;
        RECT 1026.010 10.480 1090.510 651.265 ;
        RECT 1016.110 10.240 1090.510 10.480 ;
        RECT 1092.910 10.480 1093.810 651.265 ;
        RECT 1096.210 10.480 1097.110 651.265 ;
        RECT 1099.510 10.480 1100.410 651.265 ;
        RECT 1102.810 10.480 1167.310 651.265 ;
        RECT 1092.910 10.240 1167.310 10.480 ;
        RECT 1169.710 10.480 1170.610 651.265 ;
        RECT 1173.010 10.480 1173.910 651.265 ;
        RECT 1176.310 10.480 1177.210 651.265 ;
        RECT 1179.610 10.480 1244.110 651.265 ;
        RECT 1169.710 10.240 1244.110 10.480 ;
        RECT 1246.510 10.480 1247.410 651.265 ;
        RECT 1249.810 10.480 1250.710 651.265 ;
        RECT 1253.110 10.480 1254.010 651.265 ;
        RECT 1256.410 10.480 1320.910 651.265 ;
        RECT 1246.510 10.240 1320.910 10.480 ;
        RECT 1323.310 10.480 1324.210 651.265 ;
        RECT 1326.610 10.480 1327.510 651.265 ;
        RECT 1329.910 10.480 1330.810 651.265 ;
        RECT 1333.210 10.480 1397.710 651.265 ;
        RECT 1323.310 10.240 1397.710 10.480 ;
        RECT 1400.110 10.480 1401.010 651.265 ;
        RECT 1403.410 10.480 1404.310 651.265 ;
        RECT 1406.710 10.480 1407.610 651.265 ;
        RECT 1410.010 10.480 1474.510 651.265 ;
        RECT 1400.110 10.240 1474.510 10.480 ;
        RECT 1476.910 10.480 1477.810 651.265 ;
        RECT 1480.210 10.480 1481.110 651.265 ;
        RECT 1483.510 10.480 1484.410 651.265 ;
        RECT 1486.810 10.480 1551.310 651.265 ;
        RECT 1476.910 10.240 1551.310 10.480 ;
        RECT 1553.710 10.480 1554.610 651.265 ;
        RECT 1557.010 10.480 1557.910 651.265 ;
        RECT 1560.310 10.480 1561.210 651.265 ;
        RECT 1563.610 10.480 1628.110 651.265 ;
        RECT 1553.710 10.240 1628.110 10.480 ;
        RECT 1630.510 10.480 1631.410 651.265 ;
        RECT 1633.810 10.480 1634.710 651.265 ;
        RECT 1637.110 10.480 1638.010 651.265 ;
        RECT 1640.410 10.480 1704.910 651.265 ;
        RECT 1630.510 10.240 1704.910 10.480 ;
        RECT 1707.310 10.480 1708.210 651.265 ;
        RECT 1710.610 10.480 1711.510 651.265 ;
        RECT 1713.910 10.480 1714.810 651.265 ;
        RECT 1717.210 10.480 1781.710 651.265 ;
        RECT 1707.310 10.240 1781.710 10.480 ;
        RECT 1784.110 10.480 1785.010 651.265 ;
        RECT 1787.410 10.480 1788.310 651.265 ;
        RECT 1790.710 10.480 1791.610 651.265 ;
        RECT 1794.010 10.480 1858.510 651.265 ;
        RECT 1784.110 10.240 1858.510 10.480 ;
        RECT 1860.910 10.480 1861.810 651.265 ;
        RECT 1864.210 10.480 1865.110 651.265 ;
        RECT 1867.510 10.480 1868.410 651.265 ;
        RECT 1870.810 10.480 1935.310 651.265 ;
        RECT 1860.910 10.240 1935.310 10.480 ;
        RECT 1937.710 10.480 1938.610 651.265 ;
        RECT 1941.010 10.480 1941.910 651.265 ;
        RECT 1944.310 10.480 1945.210 651.265 ;
        RECT 1947.610 10.480 2012.110 651.265 ;
        RECT 1937.710 10.240 2012.110 10.480 ;
        RECT 2014.510 10.480 2015.410 651.265 ;
        RECT 2017.810 10.480 2018.710 651.265 ;
        RECT 2021.110 10.480 2022.010 651.265 ;
        RECT 2024.410 10.480 2088.910 651.265 ;
        RECT 2014.510 10.240 2088.910 10.480 ;
        RECT 2091.310 10.480 2092.210 651.265 ;
        RECT 2094.610 10.480 2095.510 651.265 ;
        RECT 2097.910 10.480 2098.810 651.265 ;
        RECT 2101.210 10.480 2165.710 651.265 ;
        RECT 2091.310 10.240 2165.710 10.480 ;
        RECT 2168.110 10.480 2169.010 651.265 ;
        RECT 2171.410 10.480 2172.310 651.265 ;
        RECT 2174.710 10.480 2175.610 651.265 ;
        RECT 2178.010 10.480 2242.510 651.265 ;
        RECT 2168.110 10.240 2242.510 10.480 ;
        RECT 2244.910 10.480 2245.810 651.265 ;
        RECT 2248.210 10.480 2249.110 651.265 ;
        RECT 2251.510 10.480 2252.410 651.265 ;
        RECT 2254.810 10.480 2319.310 651.265 ;
        RECT 2244.910 10.240 2319.310 10.480 ;
        RECT 2321.710 10.480 2322.610 651.265 ;
        RECT 2325.010 10.480 2325.910 651.265 ;
        RECT 2328.310 10.480 2329.210 651.265 ;
        RECT 2331.610 10.480 2396.110 651.265 ;
        RECT 2321.710 10.240 2396.110 10.480 ;
        RECT 2398.510 10.480 2399.410 651.265 ;
        RECT 2401.810 10.480 2402.710 651.265 ;
        RECT 2405.110 10.480 2406.010 651.265 ;
        RECT 2408.410 10.480 2472.910 651.265 ;
        RECT 2398.510 10.240 2472.910 10.480 ;
        RECT 2475.310 10.480 2476.210 651.265 ;
        RECT 2478.610 10.480 2479.510 651.265 ;
        RECT 2481.910 10.480 2482.810 651.265 ;
        RECT 2485.210 10.480 2549.710 651.265 ;
        RECT 2475.310 10.240 2549.710 10.480 ;
        RECT 2552.110 10.480 2553.010 651.265 ;
        RECT 2555.410 10.480 2556.310 651.265 ;
        RECT 2558.710 10.480 2559.610 651.265 ;
        RECT 2562.010 10.480 2626.510 651.265 ;
        RECT 2552.110 10.240 2626.510 10.480 ;
        RECT 2628.910 10.480 2629.810 651.265 ;
        RECT 2632.210 10.480 2633.110 651.265 ;
        RECT 2635.510 10.480 2636.410 651.265 ;
        RECT 2638.810 10.480 2692.735 651.265 ;
        RECT 2628.910 10.240 2692.735 10.480 ;
        RECT 187.245 9.695 2692.735 10.240 ;
      LAYER met5 ;
        RECT 1391.810 96.100 2256.370 417.300 ;
  END
END RAM_512x64
END LIBRARY

