magic
tech sky130A
magscale 1 2
timestamp 1608837809
<< obsli1 >>
rect 1104 2159 143031 141457
<< obsm1 >>
rect 290 1232 143598 142180
<< metal2 >>
rect 386 143200 442 144000
rect 1214 143200 1270 144000
rect 2042 143200 2098 144000
rect 2870 143200 2926 144000
rect 3698 143200 3754 144000
rect 4526 143200 4582 144000
rect 5354 143200 5410 144000
rect 6182 143200 6238 144000
rect 7010 143200 7066 144000
rect 7838 143200 7894 144000
rect 8666 143200 8722 144000
rect 9494 143200 9550 144000
rect 10322 143200 10378 144000
rect 11150 143200 11206 144000
rect 11978 143200 12034 144000
rect 12806 143200 12862 144000
rect 13634 143200 13690 144000
rect 14462 143200 14518 144000
rect 15290 143200 15346 144000
rect 16118 143200 16174 144000
rect 16946 143200 17002 144000
rect 17774 143200 17830 144000
rect 18694 143200 18750 144000
rect 19522 143200 19578 144000
rect 20350 143200 20406 144000
rect 21178 143200 21234 144000
rect 22006 143200 22062 144000
rect 22834 143200 22890 144000
rect 23662 143200 23718 144000
rect 24490 143200 24546 144000
rect 25318 143200 25374 144000
rect 26146 143200 26202 144000
rect 26974 143200 27030 144000
rect 27802 143200 27858 144000
rect 28630 143200 28686 144000
rect 29458 143200 29514 144000
rect 30286 143200 30342 144000
rect 31114 143200 31170 144000
rect 31942 143200 31998 144000
rect 32770 143200 32826 144000
rect 33598 143200 33654 144000
rect 34426 143200 34482 144000
rect 35254 143200 35310 144000
rect 36082 143200 36138 144000
rect 37002 143200 37058 144000
rect 37830 143200 37886 144000
rect 38658 143200 38714 144000
rect 39486 143200 39542 144000
rect 40314 143200 40370 144000
rect 41142 143200 41198 144000
rect 41970 143200 42026 144000
rect 42798 143200 42854 144000
rect 43626 143200 43682 144000
rect 44454 143200 44510 144000
rect 45282 143200 45338 144000
rect 46110 143200 46166 144000
rect 46938 143200 46994 144000
rect 47766 143200 47822 144000
rect 48594 143200 48650 144000
rect 49422 143200 49478 144000
rect 50250 143200 50306 144000
rect 51078 143200 51134 144000
rect 51906 143200 51962 144000
rect 52734 143200 52790 144000
rect 53562 143200 53618 144000
rect 54482 143200 54538 144000
rect 55310 143200 55366 144000
rect 56138 143200 56194 144000
rect 56966 143200 57022 144000
rect 57794 143200 57850 144000
rect 58622 143200 58678 144000
rect 59450 143200 59506 144000
rect 60278 143200 60334 144000
rect 61106 143200 61162 144000
rect 61934 143200 61990 144000
rect 62762 143200 62818 144000
rect 63590 143200 63646 144000
rect 64418 143200 64474 144000
rect 65246 143200 65302 144000
rect 66074 143200 66130 144000
rect 66902 143200 66958 144000
rect 67730 143200 67786 144000
rect 68558 143200 68614 144000
rect 69386 143200 69442 144000
rect 70214 143200 70270 144000
rect 71042 143200 71098 144000
rect 71870 143200 71926 144000
rect 72790 143200 72846 144000
rect 73618 143200 73674 144000
rect 74446 143200 74502 144000
rect 75274 143200 75330 144000
rect 76102 143200 76158 144000
rect 76930 143200 76986 144000
rect 77758 143200 77814 144000
rect 78586 143200 78642 144000
rect 79414 143200 79470 144000
rect 80242 143200 80298 144000
rect 81070 143200 81126 144000
rect 81898 143200 81954 144000
rect 82726 143200 82782 144000
rect 83554 143200 83610 144000
rect 84382 143200 84438 144000
rect 85210 143200 85266 144000
rect 86038 143200 86094 144000
rect 86866 143200 86922 144000
rect 87694 143200 87750 144000
rect 88522 143200 88578 144000
rect 89350 143200 89406 144000
rect 90178 143200 90234 144000
rect 91098 143200 91154 144000
rect 91926 143200 91982 144000
rect 92754 143200 92810 144000
rect 93582 143200 93638 144000
rect 94410 143200 94466 144000
rect 95238 143200 95294 144000
rect 96066 143200 96122 144000
rect 96894 143200 96950 144000
rect 97722 143200 97778 144000
rect 98550 143200 98606 144000
rect 99378 143200 99434 144000
rect 100206 143200 100262 144000
rect 101034 143200 101090 144000
rect 101862 143200 101918 144000
rect 102690 143200 102746 144000
rect 103518 143200 103574 144000
rect 104346 143200 104402 144000
rect 105174 143200 105230 144000
rect 106002 143200 106058 144000
rect 106830 143200 106886 144000
rect 107658 143200 107714 144000
rect 108578 143200 108634 144000
rect 109406 143200 109462 144000
rect 110234 143200 110290 144000
rect 111062 143200 111118 144000
rect 111890 143200 111946 144000
rect 112718 143200 112774 144000
rect 113546 143200 113602 144000
rect 114374 143200 114430 144000
rect 115202 143200 115258 144000
rect 116030 143200 116086 144000
rect 116858 143200 116914 144000
rect 117686 143200 117742 144000
rect 118514 143200 118570 144000
rect 119342 143200 119398 144000
rect 120170 143200 120226 144000
rect 120998 143200 121054 144000
rect 121826 143200 121882 144000
rect 122654 143200 122710 144000
rect 123482 143200 123538 144000
rect 124310 143200 124366 144000
rect 125138 143200 125194 144000
rect 125966 143200 126022 144000
rect 126886 143200 126942 144000
rect 127714 143200 127770 144000
rect 128542 143200 128598 144000
rect 129370 143200 129426 144000
rect 130198 143200 130254 144000
rect 131026 143200 131082 144000
rect 131854 143200 131910 144000
rect 132682 143200 132738 144000
rect 133510 143200 133566 144000
rect 134338 143200 134394 144000
rect 135166 143200 135222 144000
rect 135994 143200 136050 144000
rect 136822 143200 136878 144000
rect 137650 143200 137706 144000
rect 138478 143200 138534 144000
rect 139306 143200 139362 144000
rect 140134 143200 140190 144000
rect 140962 143200 141018 144000
rect 141790 143200 141846 144000
rect 142618 143200 142674 144000
rect 143446 143200 143502 144000
rect 294 0 350 800
rect 938 0 994 800
rect 1582 0 1638 800
rect 2318 0 2374 800
rect 2962 0 3018 800
rect 3606 0 3662 800
rect 4342 0 4398 800
rect 4986 0 5042 800
rect 5722 0 5778 800
rect 6366 0 6422 800
rect 7010 0 7066 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9770 0 9826 800
rect 10414 0 10470 800
rect 11150 0 11206 800
rect 11794 0 11850 800
rect 12438 0 12494 800
rect 13174 0 13230 800
rect 13818 0 13874 800
rect 14554 0 14610 800
rect 15198 0 15254 800
rect 15842 0 15898 800
rect 16578 0 16634 800
rect 17222 0 17278 800
rect 17866 0 17922 800
rect 18602 0 18658 800
rect 19246 0 19302 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 22006 0 22062 800
rect 22650 0 22706 800
rect 23294 0 23350 800
rect 24030 0 24086 800
rect 24674 0 24730 800
rect 25410 0 25466 800
rect 26054 0 26110 800
rect 26698 0 26754 800
rect 27434 0 27490 800
rect 28078 0 28134 800
rect 28814 0 28870 800
rect 29458 0 29514 800
rect 30102 0 30158 800
rect 30838 0 30894 800
rect 31482 0 31538 800
rect 32126 0 32182 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34242 0 34298 800
rect 34886 0 34942 800
rect 35530 0 35586 800
rect 36266 0 36322 800
rect 36910 0 36966 800
rect 37646 0 37702 800
rect 38290 0 38346 800
rect 38934 0 38990 800
rect 39670 0 39726 800
rect 40314 0 40370 800
rect 40958 0 41014 800
rect 41694 0 41750 800
rect 42338 0 42394 800
rect 43074 0 43130 800
rect 43718 0 43774 800
rect 44362 0 44418 800
rect 45098 0 45154 800
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 47122 0 47178 800
rect 47766 0 47822 800
rect 48502 0 48558 800
rect 49146 0 49202 800
rect 49790 0 49846 800
rect 50526 0 50582 800
rect 51170 0 51226 800
rect 51906 0 51962 800
rect 52550 0 52606 800
rect 53194 0 53250 800
rect 53930 0 53986 800
rect 54574 0 54630 800
rect 55218 0 55274 800
rect 55954 0 56010 800
rect 56598 0 56654 800
rect 57334 0 57390 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59358 0 59414 800
rect 60002 0 60058 800
rect 60738 0 60794 800
rect 61382 0 61438 800
rect 62026 0 62082 800
rect 62762 0 62818 800
rect 63406 0 63462 800
rect 64050 0 64106 800
rect 64786 0 64842 800
rect 65430 0 65486 800
rect 66166 0 66222 800
rect 66810 0 66866 800
rect 67454 0 67510 800
rect 68190 0 68246 800
rect 68834 0 68890 800
rect 69478 0 69534 800
rect 70214 0 70270 800
rect 70858 0 70914 800
rect 71594 0 71650 800
rect 72238 0 72294 800
rect 72882 0 72938 800
rect 73618 0 73674 800
rect 74262 0 74318 800
rect 74998 0 75054 800
rect 75642 0 75698 800
rect 76286 0 76342 800
rect 77022 0 77078 800
rect 77666 0 77722 800
rect 78310 0 78366 800
rect 79046 0 79102 800
rect 79690 0 79746 800
rect 80426 0 80482 800
rect 81070 0 81126 800
rect 81714 0 81770 800
rect 82450 0 82506 800
rect 83094 0 83150 800
rect 83738 0 83794 800
rect 84474 0 84530 800
rect 85118 0 85174 800
rect 85854 0 85910 800
rect 86498 0 86554 800
rect 87142 0 87198 800
rect 87878 0 87934 800
rect 88522 0 88578 800
rect 89258 0 89314 800
rect 89902 0 89958 800
rect 90546 0 90602 800
rect 91282 0 91338 800
rect 91926 0 91982 800
rect 92570 0 92626 800
rect 93306 0 93362 800
rect 93950 0 94006 800
rect 94686 0 94742 800
rect 95330 0 95386 800
rect 95974 0 96030 800
rect 96710 0 96766 800
rect 97354 0 97410 800
rect 98090 0 98146 800
rect 98734 0 98790 800
rect 99378 0 99434 800
rect 100114 0 100170 800
rect 100758 0 100814 800
rect 101402 0 101458 800
rect 102138 0 102194 800
rect 102782 0 102838 800
rect 103518 0 103574 800
rect 104162 0 104218 800
rect 104806 0 104862 800
rect 105542 0 105598 800
rect 106186 0 106242 800
rect 106830 0 106886 800
rect 107566 0 107622 800
rect 108210 0 108266 800
rect 108946 0 109002 800
rect 109590 0 109646 800
rect 110234 0 110290 800
rect 110970 0 111026 800
rect 111614 0 111670 800
rect 112350 0 112406 800
rect 112994 0 113050 800
rect 113638 0 113694 800
rect 114374 0 114430 800
rect 115018 0 115074 800
rect 115662 0 115718 800
rect 116398 0 116454 800
rect 117042 0 117098 800
rect 117778 0 117834 800
rect 118422 0 118478 800
rect 119066 0 119122 800
rect 119802 0 119858 800
rect 120446 0 120502 800
rect 121182 0 121238 800
rect 121826 0 121882 800
rect 122470 0 122526 800
rect 123206 0 123262 800
rect 123850 0 123906 800
rect 124494 0 124550 800
rect 125230 0 125286 800
rect 125874 0 125930 800
rect 126610 0 126666 800
rect 127254 0 127310 800
rect 127898 0 127954 800
rect 128634 0 128690 800
rect 129278 0 129334 800
rect 129922 0 129978 800
rect 130658 0 130714 800
rect 131302 0 131358 800
rect 132038 0 132094 800
rect 132682 0 132738 800
rect 133326 0 133382 800
rect 134062 0 134118 800
rect 134706 0 134762 800
rect 135442 0 135498 800
rect 136086 0 136142 800
rect 136730 0 136786 800
rect 137466 0 137522 800
rect 138110 0 138166 800
rect 138754 0 138810 800
rect 139490 0 139546 800
rect 140134 0 140190 800
rect 140870 0 140926 800
rect 141514 0 141570 800
rect 142158 0 142214 800
rect 142894 0 142950 800
rect 143538 0 143594 800
<< obsm2 >>
rect 296 143144 330 143585
rect 498 143144 1158 143585
rect 1326 143144 1986 143585
rect 2154 143144 2814 143585
rect 2982 143144 3642 143585
rect 3810 143144 4470 143585
rect 4638 143144 5298 143585
rect 5466 143144 6126 143585
rect 6294 143144 6954 143585
rect 7122 143144 7782 143585
rect 7950 143144 8610 143585
rect 8778 143144 9438 143585
rect 9606 143144 10266 143585
rect 10434 143144 11094 143585
rect 11262 143144 11922 143585
rect 12090 143144 12750 143585
rect 12918 143144 13578 143585
rect 13746 143144 14406 143585
rect 14574 143144 15234 143585
rect 15402 143144 16062 143585
rect 16230 143144 16890 143585
rect 17058 143144 17718 143585
rect 17886 143144 18638 143585
rect 18806 143144 19466 143585
rect 19634 143144 20294 143585
rect 20462 143144 21122 143585
rect 21290 143144 21950 143585
rect 22118 143144 22778 143585
rect 22946 143144 23606 143585
rect 23774 143144 24434 143585
rect 24602 143144 25262 143585
rect 25430 143144 26090 143585
rect 26258 143144 26918 143585
rect 27086 143144 27746 143585
rect 27914 143144 28574 143585
rect 28742 143144 29402 143585
rect 29570 143144 30230 143585
rect 30398 143144 31058 143585
rect 31226 143144 31886 143585
rect 32054 143144 32714 143585
rect 32882 143144 33542 143585
rect 33710 143144 34370 143585
rect 34538 143144 35198 143585
rect 35366 143144 36026 143585
rect 36194 143144 36946 143585
rect 37114 143144 37774 143585
rect 37942 143144 38602 143585
rect 38770 143144 39430 143585
rect 39598 143144 40258 143585
rect 40426 143144 41086 143585
rect 41254 143144 41914 143585
rect 42082 143144 42742 143585
rect 42910 143144 43570 143585
rect 43738 143144 44398 143585
rect 44566 143144 45226 143585
rect 45394 143144 46054 143585
rect 46222 143144 46882 143585
rect 47050 143144 47710 143585
rect 47878 143144 48538 143585
rect 48706 143144 49366 143585
rect 49534 143144 50194 143585
rect 50362 143144 51022 143585
rect 51190 143144 51850 143585
rect 52018 143144 52678 143585
rect 52846 143144 53506 143585
rect 53674 143144 54426 143585
rect 54594 143144 55254 143585
rect 55422 143144 56082 143585
rect 56250 143144 56910 143585
rect 57078 143144 57738 143585
rect 57906 143144 58566 143585
rect 58734 143144 59394 143585
rect 59562 143144 60222 143585
rect 60390 143144 61050 143585
rect 61218 143144 61878 143585
rect 62046 143144 62706 143585
rect 62874 143144 63534 143585
rect 63702 143144 64362 143585
rect 64530 143144 65190 143585
rect 65358 143144 66018 143585
rect 66186 143144 66846 143585
rect 67014 143144 67674 143585
rect 67842 143144 68502 143585
rect 68670 143144 69330 143585
rect 69498 143144 70158 143585
rect 70326 143144 70986 143585
rect 71154 143144 71814 143585
rect 71982 143144 72734 143585
rect 72902 143144 73562 143585
rect 73730 143144 74390 143585
rect 74558 143144 75218 143585
rect 75386 143144 76046 143585
rect 76214 143144 76874 143585
rect 77042 143144 77702 143585
rect 77870 143144 78530 143585
rect 78698 143144 79358 143585
rect 79526 143144 80186 143585
rect 80354 143144 81014 143585
rect 81182 143144 81842 143585
rect 82010 143144 82670 143585
rect 82838 143144 83498 143585
rect 83666 143144 84326 143585
rect 84494 143144 85154 143585
rect 85322 143144 85982 143585
rect 86150 143144 86810 143585
rect 86978 143144 87638 143585
rect 87806 143144 88466 143585
rect 88634 143144 89294 143585
rect 89462 143144 90122 143585
rect 90290 143144 91042 143585
rect 91210 143144 91870 143585
rect 92038 143144 92698 143585
rect 92866 143144 93526 143585
rect 93694 143144 94354 143585
rect 94522 143144 95182 143585
rect 95350 143144 96010 143585
rect 96178 143144 96838 143585
rect 97006 143144 97666 143585
rect 97834 143144 98494 143585
rect 98662 143144 99322 143585
rect 99490 143144 100150 143585
rect 100318 143144 100978 143585
rect 101146 143144 101806 143585
rect 101974 143144 102634 143585
rect 102802 143144 103462 143585
rect 103630 143144 104290 143585
rect 104458 143144 105118 143585
rect 105286 143144 105946 143585
rect 106114 143144 106774 143585
rect 106942 143144 107602 143585
rect 107770 143144 108522 143585
rect 108690 143144 109350 143585
rect 109518 143144 110178 143585
rect 110346 143144 111006 143585
rect 111174 143144 111834 143585
rect 112002 143144 112662 143585
rect 112830 143144 113490 143585
rect 113658 143144 114318 143585
rect 114486 143144 115146 143585
rect 115314 143144 115974 143585
rect 116142 143144 116802 143585
rect 116970 143144 117630 143585
rect 117798 143144 118458 143585
rect 118626 143144 119286 143585
rect 119454 143144 120114 143585
rect 120282 143144 120942 143585
rect 121110 143144 121770 143585
rect 121938 143144 122598 143585
rect 122766 143144 123426 143585
rect 123594 143144 124254 143585
rect 124422 143144 125082 143585
rect 125250 143144 125910 143585
rect 126078 143144 126830 143585
rect 126998 143144 127658 143585
rect 127826 143144 128486 143585
rect 128654 143144 129314 143585
rect 129482 143144 130142 143585
rect 130310 143144 130970 143585
rect 131138 143144 131798 143585
rect 131966 143144 132626 143585
rect 132794 143144 133454 143585
rect 133622 143144 134282 143585
rect 134450 143144 135110 143585
rect 135278 143144 135938 143585
rect 136106 143144 136766 143585
rect 136934 143144 137594 143585
rect 137762 143144 138422 143585
rect 138590 143144 139250 143585
rect 139418 143144 140078 143585
rect 140246 143144 140906 143585
rect 141074 143144 141734 143585
rect 141902 143144 142562 143585
rect 142730 143144 143390 143585
rect 143558 143144 143592 143585
rect 296 856 143592 143144
rect 406 303 882 856
rect 1050 303 1526 856
rect 1694 303 2262 856
rect 2430 303 2906 856
rect 3074 303 3550 856
rect 3718 303 4286 856
rect 4454 303 4930 856
rect 5098 303 5666 856
rect 5834 303 6310 856
rect 6478 303 6954 856
rect 7122 303 7690 856
rect 7858 303 8334 856
rect 8502 303 8978 856
rect 9146 303 9714 856
rect 9882 303 10358 856
rect 10526 303 11094 856
rect 11262 303 11738 856
rect 11906 303 12382 856
rect 12550 303 13118 856
rect 13286 303 13762 856
rect 13930 303 14498 856
rect 14666 303 15142 856
rect 15310 303 15786 856
rect 15954 303 16522 856
rect 16690 303 17166 856
rect 17334 303 17810 856
rect 17978 303 18546 856
rect 18714 303 19190 856
rect 19358 303 19926 856
rect 20094 303 20570 856
rect 20738 303 21214 856
rect 21382 303 21950 856
rect 22118 303 22594 856
rect 22762 303 23238 856
rect 23406 303 23974 856
rect 24142 303 24618 856
rect 24786 303 25354 856
rect 25522 303 25998 856
rect 26166 303 26642 856
rect 26810 303 27378 856
rect 27546 303 28022 856
rect 28190 303 28758 856
rect 28926 303 29402 856
rect 29570 303 30046 856
rect 30214 303 30782 856
rect 30950 303 31426 856
rect 31594 303 32070 856
rect 32238 303 32806 856
rect 32974 303 33450 856
rect 33618 303 34186 856
rect 34354 303 34830 856
rect 34998 303 35474 856
rect 35642 303 36210 856
rect 36378 303 36854 856
rect 37022 303 37590 856
rect 37758 303 38234 856
rect 38402 303 38878 856
rect 39046 303 39614 856
rect 39782 303 40258 856
rect 40426 303 40902 856
rect 41070 303 41638 856
rect 41806 303 42282 856
rect 42450 303 43018 856
rect 43186 303 43662 856
rect 43830 303 44306 856
rect 44474 303 45042 856
rect 45210 303 45686 856
rect 45854 303 46330 856
rect 46498 303 47066 856
rect 47234 303 47710 856
rect 47878 303 48446 856
rect 48614 303 49090 856
rect 49258 303 49734 856
rect 49902 303 50470 856
rect 50638 303 51114 856
rect 51282 303 51850 856
rect 52018 303 52494 856
rect 52662 303 53138 856
rect 53306 303 53874 856
rect 54042 303 54518 856
rect 54686 303 55162 856
rect 55330 303 55898 856
rect 56066 303 56542 856
rect 56710 303 57278 856
rect 57446 303 57922 856
rect 58090 303 58566 856
rect 58734 303 59302 856
rect 59470 303 59946 856
rect 60114 303 60682 856
rect 60850 303 61326 856
rect 61494 303 61970 856
rect 62138 303 62706 856
rect 62874 303 63350 856
rect 63518 303 63994 856
rect 64162 303 64730 856
rect 64898 303 65374 856
rect 65542 303 66110 856
rect 66278 303 66754 856
rect 66922 303 67398 856
rect 67566 303 68134 856
rect 68302 303 68778 856
rect 68946 303 69422 856
rect 69590 303 70158 856
rect 70326 303 70802 856
rect 70970 303 71538 856
rect 71706 303 72182 856
rect 72350 303 72826 856
rect 72994 303 73562 856
rect 73730 303 74206 856
rect 74374 303 74942 856
rect 75110 303 75586 856
rect 75754 303 76230 856
rect 76398 303 76966 856
rect 77134 303 77610 856
rect 77778 303 78254 856
rect 78422 303 78990 856
rect 79158 303 79634 856
rect 79802 303 80370 856
rect 80538 303 81014 856
rect 81182 303 81658 856
rect 81826 303 82394 856
rect 82562 303 83038 856
rect 83206 303 83682 856
rect 83850 303 84418 856
rect 84586 303 85062 856
rect 85230 303 85798 856
rect 85966 303 86442 856
rect 86610 303 87086 856
rect 87254 303 87822 856
rect 87990 303 88466 856
rect 88634 303 89202 856
rect 89370 303 89846 856
rect 90014 303 90490 856
rect 90658 303 91226 856
rect 91394 303 91870 856
rect 92038 303 92514 856
rect 92682 303 93250 856
rect 93418 303 93894 856
rect 94062 303 94630 856
rect 94798 303 95274 856
rect 95442 303 95918 856
rect 96086 303 96654 856
rect 96822 303 97298 856
rect 97466 303 98034 856
rect 98202 303 98678 856
rect 98846 303 99322 856
rect 99490 303 100058 856
rect 100226 303 100702 856
rect 100870 303 101346 856
rect 101514 303 102082 856
rect 102250 303 102726 856
rect 102894 303 103462 856
rect 103630 303 104106 856
rect 104274 303 104750 856
rect 104918 303 105486 856
rect 105654 303 106130 856
rect 106298 303 106774 856
rect 106942 303 107510 856
rect 107678 303 108154 856
rect 108322 303 108890 856
rect 109058 303 109534 856
rect 109702 303 110178 856
rect 110346 303 110914 856
rect 111082 303 111558 856
rect 111726 303 112294 856
rect 112462 303 112938 856
rect 113106 303 113582 856
rect 113750 303 114318 856
rect 114486 303 114962 856
rect 115130 303 115606 856
rect 115774 303 116342 856
rect 116510 303 116986 856
rect 117154 303 117722 856
rect 117890 303 118366 856
rect 118534 303 119010 856
rect 119178 303 119746 856
rect 119914 303 120390 856
rect 120558 303 121126 856
rect 121294 303 121770 856
rect 121938 303 122414 856
rect 122582 303 123150 856
rect 123318 303 123794 856
rect 123962 303 124438 856
rect 124606 303 125174 856
rect 125342 303 125818 856
rect 125986 303 126554 856
rect 126722 303 127198 856
rect 127366 303 127842 856
rect 128010 303 128578 856
rect 128746 303 129222 856
rect 129390 303 129866 856
rect 130034 303 130602 856
rect 130770 303 131246 856
rect 131414 303 131982 856
rect 132150 303 132626 856
rect 132794 303 133270 856
rect 133438 303 134006 856
rect 134174 303 134650 856
rect 134818 303 135386 856
rect 135554 303 136030 856
rect 136198 303 136674 856
rect 136842 303 137410 856
rect 137578 303 138054 856
rect 138222 303 138698 856
rect 138866 303 139434 856
rect 139602 303 140078 856
rect 140246 303 140814 856
rect 140982 303 141458 856
rect 141626 303 142102 856
rect 142270 303 142838 856
rect 143006 303 143482 856
<< metal3 >>
rect 0 143488 800 143608
rect 0 142808 800 142928
rect 0 142128 800 142248
rect 0 141312 800 141432
rect 0 140632 800 140752
rect 0 139952 800 140072
rect 0 139272 800 139392
rect 0 138456 800 138576
rect 0 137776 800 137896
rect 0 137096 800 137216
rect 0 136416 800 136536
rect 0 135600 800 135720
rect 0 134920 800 135040
rect 0 134240 800 134360
rect 0 133424 800 133544
rect 0 132744 800 132864
rect 0 132064 800 132184
rect 0 131384 800 131504
rect 0 130568 800 130688
rect 0 129888 800 130008
rect 0 129208 800 129328
rect 0 128528 800 128648
rect 0 127712 800 127832
rect 0 127032 800 127152
rect 0 126352 800 126472
rect 0 125672 800 125792
rect 0 124856 800 124976
rect 0 124176 800 124296
rect 0 123496 800 123616
rect 0 122680 800 122800
rect 0 122000 800 122120
rect 0 121320 800 121440
rect 0 120640 800 120760
rect 0 119824 800 119944
rect 0 119144 800 119264
rect 0 118464 800 118584
rect 0 117784 800 117904
rect 0 116968 800 117088
rect 0 116288 800 116408
rect 0 115608 800 115728
rect 0 114792 800 114912
rect 0 114112 800 114232
rect 0 113432 800 113552
rect 0 112752 800 112872
rect 0 111936 800 112056
rect 0 111256 800 111376
rect 0 110576 800 110696
rect 0 109896 800 110016
rect 0 109080 800 109200
rect 0 108400 800 108520
rect 0 107720 800 107840
rect 0 107040 800 107160
rect 0 106224 800 106344
rect 0 105544 800 105664
rect 0 104864 800 104984
rect 0 104048 800 104168
rect 0 103368 800 103488
rect 0 102688 800 102808
rect 0 102008 800 102128
rect 0 101192 800 101312
rect 0 100512 800 100632
rect 0 99832 800 99952
rect 0 99152 800 99272
rect 0 98336 800 98456
rect 0 97656 800 97776
rect 0 96976 800 97096
rect 0 96296 800 96416
rect 0 95480 800 95600
rect 0 94800 800 94920
rect 0 94120 800 94240
rect 0 93304 800 93424
rect 0 92624 800 92744
rect 0 91944 800 92064
rect 0 91264 800 91384
rect 0 90448 800 90568
rect 0 89768 800 89888
rect 0 89088 800 89208
rect 0 88408 800 88528
rect 0 87592 800 87712
rect 0 86912 800 87032
rect 0 86232 800 86352
rect 0 85416 800 85536
rect 0 84736 800 84856
rect 0 84056 800 84176
rect 0 83376 800 83496
rect 0 82560 800 82680
rect 0 81880 800 82000
rect 0 81200 800 81320
rect 0 80520 800 80640
rect 0 79704 800 79824
rect 0 79024 800 79144
rect 0 78344 800 78464
rect 0 77664 800 77784
rect 0 76848 800 76968
rect 0 76168 800 76288
rect 0 75488 800 75608
rect 0 74672 800 74792
rect 0 73992 800 74112
rect 0 73312 800 73432
rect 0 72632 800 72752
rect 0 71816 800 71936
rect 0 71136 800 71256
rect 0 70456 800 70576
rect 0 69776 800 69896
rect 0 68960 800 69080
rect 0 68280 800 68400
rect 0 67600 800 67720
rect 0 66784 800 66904
rect 0 66104 800 66224
rect 0 65424 800 65544
rect 0 64744 800 64864
rect 0 63928 800 64048
rect 0 63248 800 63368
rect 0 62568 800 62688
rect 0 61888 800 62008
rect 0 61072 800 61192
rect 0 60392 800 60512
rect 0 59712 800 59832
rect 0 59032 800 59152
rect 0 58216 800 58336
rect 0 57536 800 57656
rect 0 56856 800 56976
rect 0 56040 800 56160
rect 0 55360 800 55480
rect 0 54680 800 54800
rect 0 54000 800 54120
rect 0 53184 800 53304
rect 0 52504 800 52624
rect 0 51824 800 51944
rect 0 51144 800 51264
rect 0 50328 800 50448
rect 0 49648 800 49768
rect 0 48968 800 49088
rect 0 48288 800 48408
rect 0 47472 800 47592
rect 0 46792 800 46912
rect 0 46112 800 46232
rect 0 45296 800 45416
rect 0 44616 800 44736
rect 0 43936 800 44056
rect 0 43256 800 43376
rect 0 42440 800 42560
rect 0 41760 800 41880
rect 0 41080 800 41200
rect 0 40400 800 40520
rect 0 39584 800 39704
rect 0 38904 800 39024
rect 0 38224 800 38344
rect 0 37408 800 37528
rect 0 36728 800 36848
rect 0 36048 800 36168
rect 0 35368 800 35488
rect 0 34552 800 34672
rect 0 33872 800 33992
rect 0 33192 800 33312
rect 0 32512 800 32632
rect 0 31696 800 31816
rect 0 31016 800 31136
rect 0 30336 800 30456
rect 0 29656 800 29776
rect 0 28840 800 28960
rect 0 28160 800 28280
rect 0 27480 800 27600
rect 0 26664 800 26784
rect 0 25984 800 26104
rect 0 25304 800 25424
rect 0 24624 800 24744
rect 0 23808 800 23928
rect 0 23128 800 23248
rect 0 22448 800 22568
rect 0 21768 800 21888
rect 0 20952 800 21072
rect 0 20272 800 20392
rect 0 19592 800 19712
rect 0 18776 800 18896
rect 0 18096 800 18216
rect 0 17416 800 17536
rect 0 16736 800 16856
rect 0 15920 800 16040
rect 0 15240 800 15360
rect 0 14560 800 14680
rect 0 13880 800 14000
rect 0 13064 800 13184
rect 0 12384 800 12504
rect 0 11704 800 11824
rect 0 11024 800 11144
rect 0 10208 800 10328
rect 0 9528 800 9648
rect 0 8848 800 8968
rect 0 8032 800 8152
rect 0 7352 800 7472
rect 0 6672 800 6792
rect 0 5992 800 6112
rect 0 5176 800 5296
rect 0 4496 800 4616
rect 0 3816 800 3936
rect 0 3136 800 3256
rect 0 2320 800 2440
rect 0 1640 800 1760
rect 0 960 800 1080
rect 0 280 800 400
<< obsm3 >>
rect 880 143408 142955 143581
rect 798 143008 142955 143408
rect 880 142728 142955 143008
rect 798 142328 142955 142728
rect 880 142048 142955 142328
rect 798 141512 142955 142048
rect 880 141232 142955 141512
rect 798 140832 142955 141232
rect 880 140552 142955 140832
rect 798 140152 142955 140552
rect 880 139872 142955 140152
rect 798 139472 142955 139872
rect 880 139192 142955 139472
rect 798 138656 142955 139192
rect 880 138376 142955 138656
rect 798 137976 142955 138376
rect 880 137696 142955 137976
rect 798 137296 142955 137696
rect 880 137016 142955 137296
rect 798 136616 142955 137016
rect 880 136336 142955 136616
rect 798 135800 142955 136336
rect 880 135520 142955 135800
rect 798 135120 142955 135520
rect 880 134840 142955 135120
rect 798 134440 142955 134840
rect 880 134160 142955 134440
rect 798 133624 142955 134160
rect 880 133344 142955 133624
rect 798 132944 142955 133344
rect 880 132664 142955 132944
rect 798 132264 142955 132664
rect 880 131984 142955 132264
rect 798 131584 142955 131984
rect 880 131304 142955 131584
rect 798 130768 142955 131304
rect 880 130488 142955 130768
rect 798 130088 142955 130488
rect 880 129808 142955 130088
rect 798 129408 142955 129808
rect 880 129128 142955 129408
rect 798 128728 142955 129128
rect 880 128448 142955 128728
rect 798 127912 142955 128448
rect 880 127632 142955 127912
rect 798 127232 142955 127632
rect 880 126952 142955 127232
rect 798 126552 142955 126952
rect 880 126272 142955 126552
rect 798 125872 142955 126272
rect 880 125592 142955 125872
rect 798 125056 142955 125592
rect 880 124776 142955 125056
rect 798 124376 142955 124776
rect 880 124096 142955 124376
rect 798 123696 142955 124096
rect 880 123416 142955 123696
rect 798 122880 142955 123416
rect 880 122600 142955 122880
rect 798 122200 142955 122600
rect 880 121920 142955 122200
rect 798 121520 142955 121920
rect 880 121240 142955 121520
rect 798 120840 142955 121240
rect 880 120560 142955 120840
rect 798 120024 142955 120560
rect 880 119744 142955 120024
rect 798 119344 142955 119744
rect 880 119064 142955 119344
rect 798 118664 142955 119064
rect 880 118384 142955 118664
rect 798 117984 142955 118384
rect 880 117704 142955 117984
rect 798 117168 142955 117704
rect 880 116888 142955 117168
rect 798 116488 142955 116888
rect 880 116208 142955 116488
rect 798 115808 142955 116208
rect 880 115528 142955 115808
rect 798 114992 142955 115528
rect 880 114712 142955 114992
rect 798 114312 142955 114712
rect 880 114032 142955 114312
rect 798 113632 142955 114032
rect 880 113352 142955 113632
rect 798 112952 142955 113352
rect 880 112672 142955 112952
rect 798 112136 142955 112672
rect 880 111856 142955 112136
rect 798 111456 142955 111856
rect 880 111176 142955 111456
rect 798 110776 142955 111176
rect 880 110496 142955 110776
rect 798 110096 142955 110496
rect 880 109816 142955 110096
rect 798 109280 142955 109816
rect 880 109000 142955 109280
rect 798 108600 142955 109000
rect 880 108320 142955 108600
rect 798 107920 142955 108320
rect 880 107640 142955 107920
rect 798 107240 142955 107640
rect 880 106960 142955 107240
rect 798 106424 142955 106960
rect 880 106144 142955 106424
rect 798 105744 142955 106144
rect 880 105464 142955 105744
rect 798 105064 142955 105464
rect 880 104784 142955 105064
rect 798 104248 142955 104784
rect 880 103968 142955 104248
rect 798 103568 142955 103968
rect 880 103288 142955 103568
rect 798 102888 142955 103288
rect 880 102608 142955 102888
rect 798 102208 142955 102608
rect 880 101928 142955 102208
rect 798 101392 142955 101928
rect 880 101112 142955 101392
rect 798 100712 142955 101112
rect 880 100432 142955 100712
rect 798 100032 142955 100432
rect 880 99752 142955 100032
rect 798 99352 142955 99752
rect 880 99072 142955 99352
rect 798 98536 142955 99072
rect 880 98256 142955 98536
rect 798 97856 142955 98256
rect 880 97576 142955 97856
rect 798 97176 142955 97576
rect 880 96896 142955 97176
rect 798 96496 142955 96896
rect 880 96216 142955 96496
rect 798 95680 142955 96216
rect 880 95400 142955 95680
rect 798 95000 142955 95400
rect 880 94720 142955 95000
rect 798 94320 142955 94720
rect 880 94040 142955 94320
rect 798 93504 142955 94040
rect 880 93224 142955 93504
rect 798 92824 142955 93224
rect 880 92544 142955 92824
rect 798 92144 142955 92544
rect 880 91864 142955 92144
rect 798 91464 142955 91864
rect 880 91184 142955 91464
rect 798 90648 142955 91184
rect 880 90368 142955 90648
rect 798 89968 142955 90368
rect 880 89688 142955 89968
rect 798 89288 142955 89688
rect 880 89008 142955 89288
rect 798 88608 142955 89008
rect 880 88328 142955 88608
rect 798 87792 142955 88328
rect 880 87512 142955 87792
rect 798 87112 142955 87512
rect 880 86832 142955 87112
rect 798 86432 142955 86832
rect 880 86152 142955 86432
rect 798 85616 142955 86152
rect 880 85336 142955 85616
rect 798 84936 142955 85336
rect 880 84656 142955 84936
rect 798 84256 142955 84656
rect 880 83976 142955 84256
rect 798 83576 142955 83976
rect 880 83296 142955 83576
rect 798 82760 142955 83296
rect 880 82480 142955 82760
rect 798 82080 142955 82480
rect 880 81800 142955 82080
rect 798 81400 142955 81800
rect 880 81120 142955 81400
rect 798 80720 142955 81120
rect 880 80440 142955 80720
rect 798 79904 142955 80440
rect 880 79624 142955 79904
rect 798 79224 142955 79624
rect 880 78944 142955 79224
rect 798 78544 142955 78944
rect 880 78264 142955 78544
rect 798 77864 142955 78264
rect 880 77584 142955 77864
rect 798 77048 142955 77584
rect 880 76768 142955 77048
rect 798 76368 142955 76768
rect 880 76088 142955 76368
rect 798 75688 142955 76088
rect 880 75408 142955 75688
rect 798 74872 142955 75408
rect 880 74592 142955 74872
rect 798 74192 142955 74592
rect 880 73912 142955 74192
rect 798 73512 142955 73912
rect 880 73232 142955 73512
rect 798 72832 142955 73232
rect 880 72552 142955 72832
rect 798 72016 142955 72552
rect 880 71736 142955 72016
rect 798 71336 142955 71736
rect 880 71056 142955 71336
rect 798 70656 142955 71056
rect 880 70376 142955 70656
rect 798 69976 142955 70376
rect 880 69696 142955 69976
rect 798 69160 142955 69696
rect 880 68880 142955 69160
rect 798 68480 142955 68880
rect 880 68200 142955 68480
rect 798 67800 142955 68200
rect 880 67520 142955 67800
rect 798 66984 142955 67520
rect 880 66704 142955 66984
rect 798 66304 142955 66704
rect 880 66024 142955 66304
rect 798 65624 142955 66024
rect 880 65344 142955 65624
rect 798 64944 142955 65344
rect 880 64664 142955 64944
rect 798 64128 142955 64664
rect 880 63848 142955 64128
rect 798 63448 142955 63848
rect 880 63168 142955 63448
rect 798 62768 142955 63168
rect 880 62488 142955 62768
rect 798 62088 142955 62488
rect 880 61808 142955 62088
rect 798 61272 142955 61808
rect 880 60992 142955 61272
rect 798 60592 142955 60992
rect 880 60312 142955 60592
rect 798 59912 142955 60312
rect 880 59632 142955 59912
rect 798 59232 142955 59632
rect 880 58952 142955 59232
rect 798 58416 142955 58952
rect 880 58136 142955 58416
rect 798 57736 142955 58136
rect 880 57456 142955 57736
rect 798 57056 142955 57456
rect 880 56776 142955 57056
rect 798 56240 142955 56776
rect 880 55960 142955 56240
rect 798 55560 142955 55960
rect 880 55280 142955 55560
rect 798 54880 142955 55280
rect 880 54600 142955 54880
rect 798 54200 142955 54600
rect 880 53920 142955 54200
rect 798 53384 142955 53920
rect 880 53104 142955 53384
rect 798 52704 142955 53104
rect 880 52424 142955 52704
rect 798 52024 142955 52424
rect 880 51744 142955 52024
rect 798 51344 142955 51744
rect 880 51064 142955 51344
rect 798 50528 142955 51064
rect 880 50248 142955 50528
rect 798 49848 142955 50248
rect 880 49568 142955 49848
rect 798 49168 142955 49568
rect 880 48888 142955 49168
rect 798 48488 142955 48888
rect 880 48208 142955 48488
rect 798 47672 142955 48208
rect 880 47392 142955 47672
rect 798 46992 142955 47392
rect 880 46712 142955 46992
rect 798 46312 142955 46712
rect 880 46032 142955 46312
rect 798 45496 142955 46032
rect 880 45216 142955 45496
rect 798 44816 142955 45216
rect 880 44536 142955 44816
rect 798 44136 142955 44536
rect 880 43856 142955 44136
rect 798 43456 142955 43856
rect 880 43176 142955 43456
rect 798 42640 142955 43176
rect 880 42360 142955 42640
rect 798 41960 142955 42360
rect 880 41680 142955 41960
rect 798 41280 142955 41680
rect 880 41000 142955 41280
rect 798 40600 142955 41000
rect 880 40320 142955 40600
rect 798 39784 142955 40320
rect 880 39504 142955 39784
rect 798 39104 142955 39504
rect 880 38824 142955 39104
rect 798 38424 142955 38824
rect 880 38144 142955 38424
rect 798 37608 142955 38144
rect 880 37328 142955 37608
rect 798 36928 142955 37328
rect 880 36648 142955 36928
rect 798 36248 142955 36648
rect 880 35968 142955 36248
rect 798 35568 142955 35968
rect 880 35288 142955 35568
rect 798 34752 142955 35288
rect 880 34472 142955 34752
rect 798 34072 142955 34472
rect 880 33792 142955 34072
rect 798 33392 142955 33792
rect 880 33112 142955 33392
rect 798 32712 142955 33112
rect 880 32432 142955 32712
rect 798 31896 142955 32432
rect 880 31616 142955 31896
rect 798 31216 142955 31616
rect 880 30936 142955 31216
rect 798 30536 142955 30936
rect 880 30256 142955 30536
rect 798 29856 142955 30256
rect 880 29576 142955 29856
rect 798 29040 142955 29576
rect 880 28760 142955 29040
rect 798 28360 142955 28760
rect 880 28080 142955 28360
rect 798 27680 142955 28080
rect 880 27400 142955 27680
rect 798 26864 142955 27400
rect 880 26584 142955 26864
rect 798 26184 142955 26584
rect 880 25904 142955 26184
rect 798 25504 142955 25904
rect 880 25224 142955 25504
rect 798 24824 142955 25224
rect 880 24544 142955 24824
rect 798 24008 142955 24544
rect 880 23728 142955 24008
rect 798 23328 142955 23728
rect 880 23048 142955 23328
rect 798 22648 142955 23048
rect 880 22368 142955 22648
rect 798 21968 142955 22368
rect 880 21688 142955 21968
rect 798 21152 142955 21688
rect 880 20872 142955 21152
rect 798 20472 142955 20872
rect 880 20192 142955 20472
rect 798 19792 142955 20192
rect 880 19512 142955 19792
rect 798 18976 142955 19512
rect 880 18696 142955 18976
rect 798 18296 142955 18696
rect 880 18016 142955 18296
rect 798 17616 142955 18016
rect 880 17336 142955 17616
rect 798 16936 142955 17336
rect 880 16656 142955 16936
rect 798 16120 142955 16656
rect 880 15840 142955 16120
rect 798 15440 142955 15840
rect 880 15160 142955 15440
rect 798 14760 142955 15160
rect 880 14480 142955 14760
rect 798 14080 142955 14480
rect 880 13800 142955 14080
rect 798 13264 142955 13800
rect 880 12984 142955 13264
rect 798 12584 142955 12984
rect 880 12304 142955 12584
rect 798 11904 142955 12304
rect 880 11624 142955 11904
rect 798 11224 142955 11624
rect 880 10944 142955 11224
rect 798 10408 142955 10944
rect 880 10128 142955 10408
rect 798 9728 142955 10128
rect 880 9448 142955 9728
rect 798 9048 142955 9448
rect 880 8768 142955 9048
rect 798 8232 142955 8768
rect 880 7952 142955 8232
rect 798 7552 142955 7952
rect 880 7272 142955 7552
rect 798 6872 142955 7272
rect 880 6592 142955 6872
rect 798 6192 142955 6592
rect 880 5912 142955 6192
rect 798 5376 142955 5912
rect 880 5096 142955 5376
rect 798 4696 142955 5096
rect 880 4416 142955 4696
rect 798 4016 142955 4416
rect 880 3736 142955 4016
rect 798 3336 142955 3736
rect 880 3056 142955 3336
rect 798 2520 142955 3056
rect 880 2240 142955 2520
rect 798 1840 142955 2240
rect 880 1560 142955 1840
rect 798 1160 142955 1560
rect 880 880 142955 1160
rect 798 480 142955 880
rect 880 307 142955 480
<< metal4 >>
rect 4208 2128 4528 141488
rect 4868 2176 5188 141440
rect 5528 2176 5848 141440
rect 6188 2176 6508 141440
rect 19568 2128 19888 141488
rect 20228 2176 20548 141440
rect 20888 2176 21208 141440
rect 21548 2176 21868 141440
rect 34928 2128 35248 141488
rect 35588 2176 35908 141440
rect 36248 2176 36568 141440
rect 36908 2176 37228 141440
rect 50288 2128 50608 141488
rect 50948 2176 51268 141440
rect 51608 2176 51928 141440
rect 52268 2176 52588 141440
rect 65648 2128 65968 141488
rect 66308 2176 66628 141440
rect 66968 2176 67288 141440
rect 67628 2176 67948 141440
rect 81008 2128 81328 141488
rect 81668 2176 81988 141440
rect 82328 2176 82648 141440
rect 82988 2176 83308 141440
rect 96368 2128 96688 141488
rect 97028 2176 97348 141440
rect 97688 2176 98008 141440
rect 98348 2176 98668 141440
rect 111728 2128 112048 141488
rect 112388 2176 112708 141440
rect 113048 2176 113368 141440
rect 113708 2176 114028 141440
rect 127088 2128 127408 141488
rect 127748 2176 128068 141440
rect 128408 2176 128728 141440
rect 129068 2176 129388 141440
<< obsm4 >>
rect 7419 141568 135733 143173
rect 7419 2619 19488 141568
rect 19968 141520 34848 141568
rect 19968 2619 20148 141520
rect 20628 2619 20808 141520
rect 21288 2619 21468 141520
rect 21948 2619 34848 141520
rect 35328 141520 50208 141568
rect 35328 2619 35508 141520
rect 35988 2619 36168 141520
rect 36648 2619 36828 141520
rect 37308 2619 50208 141520
rect 50688 141520 65568 141568
rect 50688 2619 50868 141520
rect 51348 2619 51528 141520
rect 52008 2619 52188 141520
rect 52668 2619 65568 141520
rect 66048 141520 80928 141568
rect 66048 2619 66228 141520
rect 66708 2619 66888 141520
rect 67368 2619 67548 141520
rect 68028 2619 80928 141520
rect 81408 141520 96288 141568
rect 81408 2619 81588 141520
rect 82068 2619 82248 141520
rect 82728 2619 82908 141520
rect 83388 2619 96288 141520
rect 96768 141520 111648 141568
rect 96768 2619 96948 141520
rect 97428 2619 97608 141520
rect 98088 2619 98268 141520
rect 98748 2619 111648 141520
rect 112128 141520 127008 141568
rect 112128 2619 112308 141520
rect 112788 2619 112968 141520
rect 113448 2619 113628 141520
rect 114108 2619 127008 141520
rect 127488 141520 135733 141568
rect 127488 2619 127668 141520
rect 128148 2619 128328 141520
rect 128808 2619 128988 141520
rect 129468 2619 135733 141520
<< labels >>
rlabel metal3 s 0 280 800 400 6 clk
port 1 nsew signal input
rlabel metal2 s 938 0 994 800 6 d_in[0]
port 2 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 d_in[100]
port 3 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 d_in[101]
port 4 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 d_in[102]
port 5 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 d_in[103]
port 6 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 d_in[104]
port 7 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 d_in[105]
port 8 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 d_in[106]
port 9 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 d_in[107]
port 10 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 d_in[108]
port 11 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 d_in[109]
port 12 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 d_in[10]
port 13 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 d_in[110]
port 14 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 d_in[111]
port 15 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 d_in[112]
port 16 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 d_in[113]
port 17 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 d_in[114]
port 18 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 d_in[115]
port 19 nsew signal input
rlabel metal2 s 79690 0 79746 800 6 d_in[116]
port 20 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 d_in[117]
port 21 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 d_in[118]
port 22 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 d_in[119]
port 23 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 d_in[11]
port 24 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 d_in[120]
port 25 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 d_in[121]
port 26 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 d_in[122]
port 27 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 d_in[123]
port 28 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 d_in[124]
port 29 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 d_in[125]
port 30 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 d_in[126]
port 31 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 d_in[127]
port 32 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 d_in[128]
port 33 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 d_in[129]
port 34 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 d_in[12]
port 35 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 d_in[130]
port 36 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 d_in[131]
port 37 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 d_in[132]
port 38 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 d_in[133]
port 39 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 d_in[134]
port 40 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 d_in[135]
port 41 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 d_in[136]
port 42 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 d_in[137]
port 43 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 d_in[138]
port 44 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 d_in[139]
port 45 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 d_in[13]
port 46 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 d_in[140]
port 47 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 d_in[141]
port 48 nsew signal input
rlabel metal2 s 97354 0 97410 800 6 d_in[142]
port 49 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 d_in[14]
port 50 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 d_in[15]
port 51 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 d_in[16]
port 52 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 d_in[17]
port 53 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 d_in[18]
port 54 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 d_in[19]
port 55 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 d_in[1]
port 56 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 d_in[20]
port 57 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 d_in[21]
port 58 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 d_in[22]
port 59 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 d_in[23]
port 60 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 d_in[24]
port 61 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 d_in[25]
port 62 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 d_in[26]
port 63 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 d_in[27]
port 64 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 d_in[28]
port 65 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 d_in[29]
port 66 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 d_in[2]
port 67 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 d_in[30]
port 68 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 d_in[31]
port 69 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 d_in[32]
port 70 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 d_in[33]
port 71 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 d_in[34]
port 72 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 d_in[35]
port 73 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 d_in[36]
port 74 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 d_in[37]
port 75 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 d_in[38]
port 76 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 d_in[39]
port 77 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 d_in[3]
port 78 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 d_in[40]
port 79 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 d_in[41]
port 80 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 d_in[42]
port 81 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 d_in[43]
port 82 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 d_in[44]
port 83 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 d_in[45]
port 84 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 d_in[46]
port 85 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 d_in[47]
port 86 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 d_in[48]
port 87 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 d_in[49]
port 88 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 d_in[4]
port 89 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 d_in[50]
port 90 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 d_in[51]
port 91 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 d_in[52]
port 92 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 d_in[53]
port 93 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 d_in[54]
port 94 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 d_in[55]
port 95 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 d_in[56]
port 96 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 d_in[57]
port 97 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 d_in[58]
port 98 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 d_in[59]
port 99 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 d_in[5]
port 100 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 d_in[60]
port 101 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 d_in[61]
port 102 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 d_in[62]
port 103 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 d_in[63]
port 104 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 d_in[64]
port 105 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 d_in[65]
port 106 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 d_in[66]
port 107 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 d_in[67]
port 108 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 d_in[68]
port 109 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 d_in[69]
port 110 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 d_in[6]
port 111 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 d_in[70]
port 112 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 d_in[71]
port 113 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 d_in[72]
port 114 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 d_in[73]
port 115 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 d_in[74]
port 116 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 d_in[75]
port 117 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 d_in[76]
port 118 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 d_in[77]
port 119 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 d_in[78]
port 120 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 d_in[79]
port 121 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 d_in[7]
port 122 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 d_in[80]
port 123 nsew signal input
rlabel metal2 s 55954 0 56010 800 6 d_in[81]
port 124 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 d_in[82]
port 125 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 d_in[83]
port 126 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 d_in[84]
port 127 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 d_in[85]
port 128 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 d_in[86]
port 129 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 d_in[87]
port 130 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 d_in[88]
port 131 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 d_in[89]
port 132 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 d_in[8]
port 133 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 d_in[90]
port 134 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 d_in[91]
port 135 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 d_in[92]
port 136 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 d_in[93]
port 137 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 d_in[94]
port 138 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 d_in[95]
port 139 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 d_in[96]
port 140 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 d_in[97]
port 141 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 d_in[98]
port 142 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 d_in[99]
port 143 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 d_in[9]
port 144 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 d_out[0]
port 145 nsew signal output
rlabel metal2 s 104806 0 104862 800 6 d_out[10]
port 146 nsew signal output
rlabel metal2 s 105542 0 105598 800 6 d_out[11]
port 147 nsew signal output
rlabel metal2 s 106186 0 106242 800 6 d_out[12]
port 148 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 d_out[13]
port 149 nsew signal output
rlabel metal2 s 107566 0 107622 800 6 d_out[14]
port 150 nsew signal output
rlabel metal2 s 108210 0 108266 800 6 d_out[15]
port 151 nsew signal output
rlabel metal2 s 108946 0 109002 800 6 d_out[16]
port 152 nsew signal output
rlabel metal2 s 109590 0 109646 800 6 d_out[17]
port 153 nsew signal output
rlabel metal2 s 110234 0 110290 800 6 d_out[18]
port 154 nsew signal output
rlabel metal2 s 110970 0 111026 800 6 d_out[19]
port 155 nsew signal output
rlabel metal2 s 98734 0 98790 800 6 d_out[1]
port 156 nsew signal output
rlabel metal2 s 111614 0 111670 800 6 d_out[20]
port 157 nsew signal output
rlabel metal2 s 112350 0 112406 800 6 d_out[21]
port 158 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 d_out[22]
port 159 nsew signal output
rlabel metal2 s 113638 0 113694 800 6 d_out[23]
port 160 nsew signal output
rlabel metal2 s 114374 0 114430 800 6 d_out[24]
port 161 nsew signal output
rlabel metal2 s 115018 0 115074 800 6 d_out[25]
port 162 nsew signal output
rlabel metal2 s 115662 0 115718 800 6 d_out[26]
port 163 nsew signal output
rlabel metal2 s 116398 0 116454 800 6 d_out[27]
port 164 nsew signal output
rlabel metal2 s 117042 0 117098 800 6 d_out[28]
port 165 nsew signal output
rlabel metal2 s 117778 0 117834 800 6 d_out[29]
port 166 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 d_out[2]
port 167 nsew signal output
rlabel metal2 s 118422 0 118478 800 6 d_out[30]
port 168 nsew signal output
rlabel metal2 s 119066 0 119122 800 6 d_out[31]
port 169 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 d_out[32]
port 170 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 d_out[33]
port 171 nsew signal output
rlabel metal2 s 121182 0 121238 800 6 d_out[34]
port 172 nsew signal output
rlabel metal2 s 121826 0 121882 800 6 d_out[35]
port 173 nsew signal output
rlabel metal2 s 122470 0 122526 800 6 d_out[36]
port 174 nsew signal output
rlabel metal2 s 123206 0 123262 800 6 d_out[37]
port 175 nsew signal output
rlabel metal2 s 123850 0 123906 800 6 d_out[38]
port 176 nsew signal output
rlabel metal2 s 124494 0 124550 800 6 d_out[39]
port 177 nsew signal output
rlabel metal2 s 100114 0 100170 800 6 d_out[3]
port 178 nsew signal output
rlabel metal2 s 125230 0 125286 800 6 d_out[40]
port 179 nsew signal output
rlabel metal2 s 125874 0 125930 800 6 d_out[41]
port 180 nsew signal output
rlabel metal2 s 126610 0 126666 800 6 d_out[42]
port 181 nsew signal output
rlabel metal2 s 127254 0 127310 800 6 d_out[43]
port 182 nsew signal output
rlabel metal2 s 127898 0 127954 800 6 d_out[44]
port 183 nsew signal output
rlabel metal2 s 128634 0 128690 800 6 d_out[45]
port 184 nsew signal output
rlabel metal2 s 129278 0 129334 800 6 d_out[46]
port 185 nsew signal output
rlabel metal2 s 129922 0 129978 800 6 d_out[47]
port 186 nsew signal output
rlabel metal2 s 130658 0 130714 800 6 d_out[48]
port 187 nsew signal output
rlabel metal2 s 131302 0 131358 800 6 d_out[49]
port 188 nsew signal output
rlabel metal2 s 100758 0 100814 800 6 d_out[4]
port 189 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 d_out[50]
port 190 nsew signal output
rlabel metal2 s 132682 0 132738 800 6 d_out[51]
port 191 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 d_out[52]
port 192 nsew signal output
rlabel metal2 s 134062 0 134118 800 6 d_out[53]
port 193 nsew signal output
rlabel metal2 s 134706 0 134762 800 6 d_out[54]
port 194 nsew signal output
rlabel metal2 s 135442 0 135498 800 6 d_out[55]
port 195 nsew signal output
rlabel metal2 s 136086 0 136142 800 6 d_out[56]
port 196 nsew signal output
rlabel metal2 s 136730 0 136786 800 6 d_out[57]
port 197 nsew signal output
rlabel metal2 s 137466 0 137522 800 6 d_out[58]
port 198 nsew signal output
rlabel metal2 s 138110 0 138166 800 6 d_out[59]
port 199 nsew signal output
rlabel metal2 s 101402 0 101458 800 6 d_out[5]
port 200 nsew signal output
rlabel metal2 s 138754 0 138810 800 6 d_out[60]
port 201 nsew signal output
rlabel metal2 s 139490 0 139546 800 6 d_out[61]
port 202 nsew signal output
rlabel metal2 s 140134 0 140190 800 6 d_out[62]
port 203 nsew signal output
rlabel metal2 s 140870 0 140926 800 6 d_out[63]
port 204 nsew signal output
rlabel metal2 s 141514 0 141570 800 6 d_out[64]
port 205 nsew signal output
rlabel metal2 s 142158 0 142214 800 6 d_out[65]
port 206 nsew signal output
rlabel metal2 s 142894 0 142950 800 6 d_out[66]
port 207 nsew signal output
rlabel metal2 s 143538 0 143594 800 6 d_out[67]
port 208 nsew signal output
rlabel metal2 s 102138 0 102194 800 6 d_out[6]
port 209 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 d_out[7]
port 210 nsew signal output
rlabel metal2 s 103518 0 103574 800 6 d_out[8]
port 211 nsew signal output
rlabel metal2 s 104162 0 104218 800 6 d_out[9]
port 212 nsew signal output
rlabel metal3 s 0 1640 800 1760 6 m_in[0]
port 213 nsew signal input
rlabel metal3 s 0 73312 800 73432 6 m_in[100]
port 214 nsew signal input
rlabel metal3 s 0 73992 800 74112 6 m_in[101]
port 215 nsew signal input
rlabel metal3 s 0 74672 800 74792 6 m_in[102]
port 216 nsew signal input
rlabel metal3 s 0 75488 800 75608 6 m_in[103]
port 217 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 m_in[104]
port 218 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 m_in[105]
port 219 nsew signal input
rlabel metal3 s 0 77664 800 77784 6 m_in[106]
port 220 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 m_in[107]
port 221 nsew signal input
rlabel metal3 s 0 79024 800 79144 6 m_in[108]
port 222 nsew signal input
rlabel metal3 s 0 79704 800 79824 6 m_in[109]
port 223 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 m_in[10]
port 224 nsew signal input
rlabel metal3 s 0 80520 800 80640 6 m_in[110]
port 225 nsew signal input
rlabel metal3 s 0 81200 800 81320 6 m_in[111]
port 226 nsew signal input
rlabel metal3 s 0 81880 800 82000 6 m_in[112]
port 227 nsew signal input
rlabel metal3 s 0 82560 800 82680 6 m_in[113]
port 228 nsew signal input
rlabel metal3 s 0 83376 800 83496 6 m_in[114]
port 229 nsew signal input
rlabel metal3 s 0 84056 800 84176 6 m_in[115]
port 230 nsew signal input
rlabel metal3 s 0 84736 800 84856 6 m_in[116]
port 231 nsew signal input
rlabel metal3 s 0 85416 800 85536 6 m_in[117]
port 232 nsew signal input
rlabel metal3 s 0 86232 800 86352 6 m_in[118]
port 233 nsew signal input
rlabel metal3 s 0 86912 800 87032 6 m_in[119]
port 234 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 m_in[11]
port 235 nsew signal input
rlabel metal3 s 0 87592 800 87712 6 m_in[120]
port 236 nsew signal input
rlabel metal3 s 0 88408 800 88528 6 m_in[121]
port 237 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 m_in[122]
port 238 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 m_in[123]
port 239 nsew signal input
rlabel metal3 s 0 90448 800 90568 6 m_in[124]
port 240 nsew signal input
rlabel metal3 s 0 91264 800 91384 6 m_in[125]
port 241 nsew signal input
rlabel metal3 s 0 91944 800 92064 6 m_in[126]
port 242 nsew signal input
rlabel metal3 s 0 92624 800 92744 6 m_in[127]
port 243 nsew signal input
rlabel metal3 s 0 93304 800 93424 6 m_in[128]
port 244 nsew signal input
rlabel metal3 s 0 94120 800 94240 6 m_in[129]
port 245 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 m_in[12]
port 246 nsew signal input
rlabel metal3 s 0 94800 800 94920 6 m_in[130]
port 247 nsew signal input
rlabel metal3 s 0 95480 800 95600 6 m_in[131]
port 248 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 m_in[13]
port 249 nsew signal input
rlabel metal3 s 0 11704 800 11824 6 m_in[14]
port 250 nsew signal input
rlabel metal3 s 0 12384 800 12504 6 m_in[15]
port 251 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 m_in[16]
port 252 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 m_in[17]
port 253 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 m_in[18]
port 254 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 m_in[19]
port 255 nsew signal input
rlabel metal3 s 0 2320 800 2440 6 m_in[1]
port 256 nsew signal input
rlabel metal3 s 0 15920 800 16040 6 m_in[20]
port 257 nsew signal input
rlabel metal3 s 0 16736 800 16856 6 m_in[21]
port 258 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 m_in[22]
port 259 nsew signal input
rlabel metal3 s 0 18096 800 18216 6 m_in[23]
port 260 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 m_in[24]
port 261 nsew signal input
rlabel metal3 s 0 19592 800 19712 6 m_in[25]
port 262 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 m_in[26]
port 263 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 m_in[27]
port 264 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 m_in[28]
port 265 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 m_in[29]
port 266 nsew signal input
rlabel metal3 s 0 3136 800 3256 6 m_in[2]
port 267 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 m_in[30]
port 268 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 m_in[31]
port 269 nsew signal input
rlabel metal3 s 0 24624 800 24744 6 m_in[32]
port 270 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 m_in[33]
port 271 nsew signal input
rlabel metal3 s 0 25984 800 26104 6 m_in[34]
port 272 nsew signal input
rlabel metal3 s 0 26664 800 26784 6 m_in[35]
port 273 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 m_in[36]
port 274 nsew signal input
rlabel metal3 s 0 28160 800 28280 6 m_in[37]
port 275 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 m_in[38]
port 276 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 m_in[39]
port 277 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 m_in[3]
port 278 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 m_in[40]
port 279 nsew signal input
rlabel metal3 s 0 31016 800 31136 6 m_in[41]
port 280 nsew signal input
rlabel metal3 s 0 31696 800 31816 6 m_in[42]
port 281 nsew signal input
rlabel metal3 s 0 32512 800 32632 6 m_in[43]
port 282 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 m_in[44]
port 283 nsew signal input
rlabel metal3 s 0 33872 800 33992 6 m_in[45]
port 284 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 m_in[46]
port 285 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 m_in[47]
port 286 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 m_in[48]
port 287 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 m_in[49]
port 288 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 m_in[4]
port 289 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 m_in[50]
port 290 nsew signal input
rlabel metal3 s 0 38224 800 38344 6 m_in[51]
port 291 nsew signal input
rlabel metal3 s 0 38904 800 39024 6 m_in[52]
port 292 nsew signal input
rlabel metal3 s 0 39584 800 39704 6 m_in[53]
port 293 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 m_in[54]
port 294 nsew signal input
rlabel metal3 s 0 41080 800 41200 6 m_in[55]
port 295 nsew signal input
rlabel metal3 s 0 41760 800 41880 6 m_in[56]
port 296 nsew signal input
rlabel metal3 s 0 42440 800 42560 6 m_in[57]
port 297 nsew signal input
rlabel metal3 s 0 43256 800 43376 6 m_in[58]
port 298 nsew signal input
rlabel metal3 s 0 43936 800 44056 6 m_in[59]
port 299 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 m_in[5]
port 300 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 m_in[60]
port 301 nsew signal input
rlabel metal3 s 0 45296 800 45416 6 m_in[61]
port 302 nsew signal input
rlabel metal3 s 0 46112 800 46232 6 m_in[62]
port 303 nsew signal input
rlabel metal3 s 0 46792 800 46912 6 m_in[63]
port 304 nsew signal input
rlabel metal3 s 0 47472 800 47592 6 m_in[64]
port 305 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 m_in[65]
port 306 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 m_in[66]
port 307 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 m_in[67]
port 308 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 m_in[68]
port 309 nsew signal input
rlabel metal3 s 0 51144 800 51264 6 m_in[69]
port 310 nsew signal input
rlabel metal3 s 0 5992 800 6112 6 m_in[6]
port 311 nsew signal input
rlabel metal3 s 0 51824 800 51944 6 m_in[70]
port 312 nsew signal input
rlabel metal3 s 0 52504 800 52624 6 m_in[71]
port 313 nsew signal input
rlabel metal3 s 0 53184 800 53304 6 m_in[72]
port 314 nsew signal input
rlabel metal3 s 0 54000 800 54120 6 m_in[73]
port 315 nsew signal input
rlabel metal3 s 0 54680 800 54800 6 m_in[74]
port 316 nsew signal input
rlabel metal3 s 0 55360 800 55480 6 m_in[75]
port 317 nsew signal input
rlabel metal3 s 0 56040 800 56160 6 m_in[76]
port 318 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 m_in[77]
port 319 nsew signal input
rlabel metal3 s 0 57536 800 57656 6 m_in[78]
port 320 nsew signal input
rlabel metal3 s 0 58216 800 58336 6 m_in[79]
port 321 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 m_in[7]
port 322 nsew signal input
rlabel metal3 s 0 59032 800 59152 6 m_in[80]
port 323 nsew signal input
rlabel metal3 s 0 59712 800 59832 6 m_in[81]
port 324 nsew signal input
rlabel metal3 s 0 60392 800 60512 6 m_in[82]
port 325 nsew signal input
rlabel metal3 s 0 61072 800 61192 6 m_in[83]
port 326 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 m_in[84]
port 327 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 m_in[85]
port 328 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 m_in[86]
port 329 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 m_in[87]
port 330 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 m_in[88]
port 331 nsew signal input
rlabel metal3 s 0 65424 800 65544 6 m_in[89]
port 332 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 m_in[8]
port 333 nsew signal input
rlabel metal3 s 0 66104 800 66224 6 m_in[90]
port 334 nsew signal input
rlabel metal3 s 0 66784 800 66904 6 m_in[91]
port 335 nsew signal input
rlabel metal3 s 0 67600 800 67720 6 m_in[92]
port 336 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 m_in[93]
port 337 nsew signal input
rlabel metal3 s 0 68960 800 69080 6 m_in[94]
port 338 nsew signal input
rlabel metal3 s 0 69776 800 69896 6 m_in[95]
port 339 nsew signal input
rlabel metal3 s 0 70456 800 70576 6 m_in[96]
port 340 nsew signal input
rlabel metal3 s 0 71136 800 71256 6 m_in[97]
port 341 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 m_in[98]
port 342 nsew signal input
rlabel metal3 s 0 72632 800 72752 6 m_in[99]
port 343 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 m_in[9]
port 344 nsew signal input
rlabel metal3 s 0 96296 800 96416 6 m_out[0]
port 345 nsew signal output
rlabel metal3 s 0 103368 800 103488 6 m_out[10]
port 346 nsew signal output
rlabel metal3 s 0 104048 800 104168 6 m_out[11]
port 347 nsew signal output
rlabel metal3 s 0 104864 800 104984 6 m_out[12]
port 348 nsew signal output
rlabel metal3 s 0 105544 800 105664 6 m_out[13]
port 349 nsew signal output
rlabel metal3 s 0 106224 800 106344 6 m_out[14]
port 350 nsew signal output
rlabel metal3 s 0 107040 800 107160 6 m_out[15]
port 351 nsew signal output
rlabel metal3 s 0 107720 800 107840 6 m_out[16]
port 352 nsew signal output
rlabel metal3 s 0 108400 800 108520 6 m_out[17]
port 353 nsew signal output
rlabel metal3 s 0 109080 800 109200 6 m_out[18]
port 354 nsew signal output
rlabel metal3 s 0 109896 800 110016 6 m_out[19]
port 355 nsew signal output
rlabel metal3 s 0 96976 800 97096 6 m_out[1]
port 356 nsew signal output
rlabel metal3 s 0 110576 800 110696 6 m_out[20]
port 357 nsew signal output
rlabel metal3 s 0 111256 800 111376 6 m_out[21]
port 358 nsew signal output
rlabel metal3 s 0 111936 800 112056 6 m_out[22]
port 359 nsew signal output
rlabel metal3 s 0 112752 800 112872 6 m_out[23]
port 360 nsew signal output
rlabel metal3 s 0 113432 800 113552 6 m_out[24]
port 361 nsew signal output
rlabel metal3 s 0 114112 800 114232 6 m_out[25]
port 362 nsew signal output
rlabel metal3 s 0 114792 800 114912 6 m_out[26]
port 363 nsew signal output
rlabel metal3 s 0 115608 800 115728 6 m_out[27]
port 364 nsew signal output
rlabel metal3 s 0 116288 800 116408 6 m_out[28]
port 365 nsew signal output
rlabel metal3 s 0 116968 800 117088 6 m_out[29]
port 366 nsew signal output
rlabel metal3 s 0 97656 800 97776 6 m_out[2]
port 367 nsew signal output
rlabel metal3 s 0 117784 800 117904 6 m_out[30]
port 368 nsew signal output
rlabel metal3 s 0 118464 800 118584 6 m_out[31]
port 369 nsew signal output
rlabel metal3 s 0 119144 800 119264 6 m_out[32]
port 370 nsew signal output
rlabel metal3 s 0 119824 800 119944 6 m_out[33]
port 371 nsew signal output
rlabel metal3 s 0 120640 800 120760 6 m_out[34]
port 372 nsew signal output
rlabel metal3 s 0 121320 800 121440 6 m_out[35]
port 373 nsew signal output
rlabel metal3 s 0 122000 800 122120 6 m_out[36]
port 374 nsew signal output
rlabel metal3 s 0 122680 800 122800 6 m_out[37]
port 375 nsew signal output
rlabel metal3 s 0 123496 800 123616 6 m_out[38]
port 376 nsew signal output
rlabel metal3 s 0 124176 800 124296 6 m_out[39]
port 377 nsew signal output
rlabel metal3 s 0 98336 800 98456 6 m_out[3]
port 378 nsew signal output
rlabel metal3 s 0 124856 800 124976 6 m_out[40]
port 379 nsew signal output
rlabel metal3 s 0 125672 800 125792 6 m_out[41]
port 380 nsew signal output
rlabel metal3 s 0 126352 800 126472 6 m_out[42]
port 381 nsew signal output
rlabel metal3 s 0 127032 800 127152 6 m_out[43]
port 382 nsew signal output
rlabel metal3 s 0 127712 800 127832 6 m_out[44]
port 383 nsew signal output
rlabel metal3 s 0 128528 800 128648 6 m_out[45]
port 384 nsew signal output
rlabel metal3 s 0 129208 800 129328 6 m_out[46]
port 385 nsew signal output
rlabel metal3 s 0 129888 800 130008 6 m_out[47]
port 386 nsew signal output
rlabel metal3 s 0 130568 800 130688 6 m_out[48]
port 387 nsew signal output
rlabel metal3 s 0 131384 800 131504 6 m_out[49]
port 388 nsew signal output
rlabel metal3 s 0 99152 800 99272 6 m_out[4]
port 389 nsew signal output
rlabel metal3 s 0 132064 800 132184 6 m_out[50]
port 390 nsew signal output
rlabel metal3 s 0 132744 800 132864 6 m_out[51]
port 391 nsew signal output
rlabel metal3 s 0 133424 800 133544 6 m_out[52]
port 392 nsew signal output
rlabel metal3 s 0 134240 800 134360 6 m_out[53]
port 393 nsew signal output
rlabel metal3 s 0 134920 800 135040 6 m_out[54]
port 394 nsew signal output
rlabel metal3 s 0 135600 800 135720 6 m_out[55]
port 395 nsew signal output
rlabel metal3 s 0 136416 800 136536 6 m_out[56]
port 396 nsew signal output
rlabel metal3 s 0 137096 800 137216 6 m_out[57]
port 397 nsew signal output
rlabel metal3 s 0 137776 800 137896 6 m_out[58]
port 398 nsew signal output
rlabel metal3 s 0 138456 800 138576 6 m_out[59]
port 399 nsew signal output
rlabel metal3 s 0 99832 800 99952 6 m_out[5]
port 400 nsew signal output
rlabel metal3 s 0 139272 800 139392 6 m_out[60]
port 401 nsew signal output
rlabel metal3 s 0 139952 800 140072 6 m_out[61]
port 402 nsew signal output
rlabel metal3 s 0 140632 800 140752 6 m_out[62]
port 403 nsew signal output
rlabel metal3 s 0 141312 800 141432 6 m_out[63]
port 404 nsew signal output
rlabel metal3 s 0 142128 800 142248 6 m_out[64]
port 405 nsew signal output
rlabel metal3 s 0 142808 800 142928 6 m_out[65]
port 406 nsew signal output
rlabel metal3 s 0 143488 800 143608 6 m_out[66]
port 407 nsew signal output
rlabel metal3 s 0 100512 800 100632 6 m_out[6]
port 408 nsew signal output
rlabel metal3 s 0 101192 800 101312 6 m_out[7]
port 409 nsew signal output
rlabel metal3 s 0 102008 800 102128 6 m_out[8]
port 410 nsew signal output
rlabel metal3 s 0 102688 800 102808 6 m_out[9]
port 411 nsew signal output
rlabel metal3 s 0 960 800 1080 6 rst
port 412 nsew signal input
rlabel metal2 s 294 0 350 800 6 stall_out
port 413 nsew signal output
rlabel metal2 s 386 143200 442 144000 6 wishbone_in[0]
port 414 nsew signal input
rlabel metal2 s 8666 143200 8722 144000 6 wishbone_in[10]
port 415 nsew signal input
rlabel metal2 s 9494 143200 9550 144000 6 wishbone_in[11]
port 416 nsew signal input
rlabel metal2 s 10322 143200 10378 144000 6 wishbone_in[12]
port 417 nsew signal input
rlabel metal2 s 11150 143200 11206 144000 6 wishbone_in[13]
port 418 nsew signal input
rlabel metal2 s 11978 143200 12034 144000 6 wishbone_in[14]
port 419 nsew signal input
rlabel metal2 s 12806 143200 12862 144000 6 wishbone_in[15]
port 420 nsew signal input
rlabel metal2 s 13634 143200 13690 144000 6 wishbone_in[16]
port 421 nsew signal input
rlabel metal2 s 14462 143200 14518 144000 6 wishbone_in[17]
port 422 nsew signal input
rlabel metal2 s 15290 143200 15346 144000 6 wishbone_in[18]
port 423 nsew signal input
rlabel metal2 s 16118 143200 16174 144000 6 wishbone_in[19]
port 424 nsew signal input
rlabel metal2 s 1214 143200 1270 144000 6 wishbone_in[1]
port 425 nsew signal input
rlabel metal2 s 16946 143200 17002 144000 6 wishbone_in[20]
port 426 nsew signal input
rlabel metal2 s 17774 143200 17830 144000 6 wishbone_in[21]
port 427 nsew signal input
rlabel metal2 s 18694 143200 18750 144000 6 wishbone_in[22]
port 428 nsew signal input
rlabel metal2 s 19522 143200 19578 144000 6 wishbone_in[23]
port 429 nsew signal input
rlabel metal2 s 20350 143200 20406 144000 6 wishbone_in[24]
port 430 nsew signal input
rlabel metal2 s 21178 143200 21234 144000 6 wishbone_in[25]
port 431 nsew signal input
rlabel metal2 s 22006 143200 22062 144000 6 wishbone_in[26]
port 432 nsew signal input
rlabel metal2 s 22834 143200 22890 144000 6 wishbone_in[27]
port 433 nsew signal input
rlabel metal2 s 23662 143200 23718 144000 6 wishbone_in[28]
port 434 nsew signal input
rlabel metal2 s 24490 143200 24546 144000 6 wishbone_in[29]
port 435 nsew signal input
rlabel metal2 s 2042 143200 2098 144000 6 wishbone_in[2]
port 436 nsew signal input
rlabel metal2 s 25318 143200 25374 144000 6 wishbone_in[30]
port 437 nsew signal input
rlabel metal2 s 26146 143200 26202 144000 6 wishbone_in[31]
port 438 nsew signal input
rlabel metal2 s 26974 143200 27030 144000 6 wishbone_in[32]
port 439 nsew signal input
rlabel metal2 s 27802 143200 27858 144000 6 wishbone_in[33]
port 440 nsew signal input
rlabel metal2 s 28630 143200 28686 144000 6 wishbone_in[34]
port 441 nsew signal input
rlabel metal2 s 29458 143200 29514 144000 6 wishbone_in[35]
port 442 nsew signal input
rlabel metal2 s 30286 143200 30342 144000 6 wishbone_in[36]
port 443 nsew signal input
rlabel metal2 s 31114 143200 31170 144000 6 wishbone_in[37]
port 444 nsew signal input
rlabel metal2 s 31942 143200 31998 144000 6 wishbone_in[38]
port 445 nsew signal input
rlabel metal2 s 32770 143200 32826 144000 6 wishbone_in[39]
port 446 nsew signal input
rlabel metal2 s 2870 143200 2926 144000 6 wishbone_in[3]
port 447 nsew signal input
rlabel metal2 s 33598 143200 33654 144000 6 wishbone_in[40]
port 448 nsew signal input
rlabel metal2 s 34426 143200 34482 144000 6 wishbone_in[41]
port 449 nsew signal input
rlabel metal2 s 35254 143200 35310 144000 6 wishbone_in[42]
port 450 nsew signal input
rlabel metal2 s 36082 143200 36138 144000 6 wishbone_in[43]
port 451 nsew signal input
rlabel metal2 s 37002 143200 37058 144000 6 wishbone_in[44]
port 452 nsew signal input
rlabel metal2 s 37830 143200 37886 144000 6 wishbone_in[45]
port 453 nsew signal input
rlabel metal2 s 38658 143200 38714 144000 6 wishbone_in[46]
port 454 nsew signal input
rlabel metal2 s 39486 143200 39542 144000 6 wishbone_in[47]
port 455 nsew signal input
rlabel metal2 s 40314 143200 40370 144000 6 wishbone_in[48]
port 456 nsew signal input
rlabel metal2 s 41142 143200 41198 144000 6 wishbone_in[49]
port 457 nsew signal input
rlabel metal2 s 3698 143200 3754 144000 6 wishbone_in[4]
port 458 nsew signal input
rlabel metal2 s 41970 143200 42026 144000 6 wishbone_in[50]
port 459 nsew signal input
rlabel metal2 s 42798 143200 42854 144000 6 wishbone_in[51]
port 460 nsew signal input
rlabel metal2 s 43626 143200 43682 144000 6 wishbone_in[52]
port 461 nsew signal input
rlabel metal2 s 44454 143200 44510 144000 6 wishbone_in[53]
port 462 nsew signal input
rlabel metal2 s 45282 143200 45338 144000 6 wishbone_in[54]
port 463 nsew signal input
rlabel metal2 s 46110 143200 46166 144000 6 wishbone_in[55]
port 464 nsew signal input
rlabel metal2 s 46938 143200 46994 144000 6 wishbone_in[56]
port 465 nsew signal input
rlabel metal2 s 47766 143200 47822 144000 6 wishbone_in[57]
port 466 nsew signal input
rlabel metal2 s 48594 143200 48650 144000 6 wishbone_in[58]
port 467 nsew signal input
rlabel metal2 s 49422 143200 49478 144000 6 wishbone_in[59]
port 468 nsew signal input
rlabel metal2 s 4526 143200 4582 144000 6 wishbone_in[5]
port 469 nsew signal input
rlabel metal2 s 50250 143200 50306 144000 6 wishbone_in[60]
port 470 nsew signal input
rlabel metal2 s 51078 143200 51134 144000 6 wishbone_in[61]
port 471 nsew signal input
rlabel metal2 s 51906 143200 51962 144000 6 wishbone_in[62]
port 472 nsew signal input
rlabel metal2 s 52734 143200 52790 144000 6 wishbone_in[63]
port 473 nsew signal input
rlabel metal2 s 53562 143200 53618 144000 6 wishbone_in[64]
port 474 nsew signal input
rlabel metal2 s 54482 143200 54538 144000 6 wishbone_in[65]
port 475 nsew signal input
rlabel metal2 s 5354 143200 5410 144000 6 wishbone_in[6]
port 476 nsew signal input
rlabel metal2 s 6182 143200 6238 144000 6 wishbone_in[7]
port 477 nsew signal input
rlabel metal2 s 7010 143200 7066 144000 6 wishbone_in[8]
port 478 nsew signal input
rlabel metal2 s 7838 143200 7894 144000 6 wishbone_in[9]
port 479 nsew signal input
rlabel metal2 s 55310 143200 55366 144000 6 wishbone_out[0]
port 480 nsew signal output
rlabel metal2 s 138478 143200 138534 144000 6 wishbone_out[100]
port 481 nsew signal output
rlabel metal2 s 139306 143200 139362 144000 6 wishbone_out[101]
port 482 nsew signal output
rlabel metal2 s 140134 143200 140190 144000 6 wishbone_out[102]
port 483 nsew signal output
rlabel metal2 s 140962 143200 141018 144000 6 wishbone_out[103]
port 484 nsew signal output
rlabel metal2 s 141790 143200 141846 144000 6 wishbone_out[104]
port 485 nsew signal output
rlabel metal2 s 142618 143200 142674 144000 6 wishbone_out[105]
port 486 nsew signal output
rlabel metal2 s 143446 143200 143502 144000 6 wishbone_out[106]
port 487 nsew signal output
rlabel metal2 s 63590 143200 63646 144000 6 wishbone_out[10]
port 488 nsew signal output
rlabel metal2 s 64418 143200 64474 144000 6 wishbone_out[11]
port 489 nsew signal output
rlabel metal2 s 65246 143200 65302 144000 6 wishbone_out[12]
port 490 nsew signal output
rlabel metal2 s 66074 143200 66130 144000 6 wishbone_out[13]
port 491 nsew signal output
rlabel metal2 s 66902 143200 66958 144000 6 wishbone_out[14]
port 492 nsew signal output
rlabel metal2 s 67730 143200 67786 144000 6 wishbone_out[15]
port 493 nsew signal output
rlabel metal2 s 68558 143200 68614 144000 6 wishbone_out[16]
port 494 nsew signal output
rlabel metal2 s 69386 143200 69442 144000 6 wishbone_out[17]
port 495 nsew signal output
rlabel metal2 s 70214 143200 70270 144000 6 wishbone_out[18]
port 496 nsew signal output
rlabel metal2 s 71042 143200 71098 144000 6 wishbone_out[19]
port 497 nsew signal output
rlabel metal2 s 56138 143200 56194 144000 6 wishbone_out[1]
port 498 nsew signal output
rlabel metal2 s 71870 143200 71926 144000 6 wishbone_out[20]
port 499 nsew signal output
rlabel metal2 s 72790 143200 72846 144000 6 wishbone_out[21]
port 500 nsew signal output
rlabel metal2 s 73618 143200 73674 144000 6 wishbone_out[22]
port 501 nsew signal output
rlabel metal2 s 74446 143200 74502 144000 6 wishbone_out[23]
port 502 nsew signal output
rlabel metal2 s 75274 143200 75330 144000 6 wishbone_out[24]
port 503 nsew signal output
rlabel metal2 s 76102 143200 76158 144000 6 wishbone_out[25]
port 504 nsew signal output
rlabel metal2 s 76930 143200 76986 144000 6 wishbone_out[26]
port 505 nsew signal output
rlabel metal2 s 77758 143200 77814 144000 6 wishbone_out[27]
port 506 nsew signal output
rlabel metal2 s 78586 143200 78642 144000 6 wishbone_out[28]
port 507 nsew signal output
rlabel metal2 s 79414 143200 79470 144000 6 wishbone_out[29]
port 508 nsew signal output
rlabel metal2 s 56966 143200 57022 144000 6 wishbone_out[2]
port 509 nsew signal output
rlabel metal2 s 80242 143200 80298 144000 6 wishbone_out[30]
port 510 nsew signal output
rlabel metal2 s 81070 143200 81126 144000 6 wishbone_out[31]
port 511 nsew signal output
rlabel metal2 s 81898 143200 81954 144000 6 wishbone_out[32]
port 512 nsew signal output
rlabel metal2 s 82726 143200 82782 144000 6 wishbone_out[33]
port 513 nsew signal output
rlabel metal2 s 83554 143200 83610 144000 6 wishbone_out[34]
port 514 nsew signal output
rlabel metal2 s 84382 143200 84438 144000 6 wishbone_out[35]
port 515 nsew signal output
rlabel metal2 s 85210 143200 85266 144000 6 wishbone_out[36]
port 516 nsew signal output
rlabel metal2 s 86038 143200 86094 144000 6 wishbone_out[37]
port 517 nsew signal output
rlabel metal2 s 86866 143200 86922 144000 6 wishbone_out[38]
port 518 nsew signal output
rlabel metal2 s 87694 143200 87750 144000 6 wishbone_out[39]
port 519 nsew signal output
rlabel metal2 s 57794 143200 57850 144000 6 wishbone_out[3]
port 520 nsew signal output
rlabel metal2 s 88522 143200 88578 144000 6 wishbone_out[40]
port 521 nsew signal output
rlabel metal2 s 89350 143200 89406 144000 6 wishbone_out[41]
port 522 nsew signal output
rlabel metal2 s 90178 143200 90234 144000 6 wishbone_out[42]
port 523 nsew signal output
rlabel metal2 s 91098 143200 91154 144000 6 wishbone_out[43]
port 524 nsew signal output
rlabel metal2 s 91926 143200 91982 144000 6 wishbone_out[44]
port 525 nsew signal output
rlabel metal2 s 92754 143200 92810 144000 6 wishbone_out[45]
port 526 nsew signal output
rlabel metal2 s 93582 143200 93638 144000 6 wishbone_out[46]
port 527 nsew signal output
rlabel metal2 s 94410 143200 94466 144000 6 wishbone_out[47]
port 528 nsew signal output
rlabel metal2 s 95238 143200 95294 144000 6 wishbone_out[48]
port 529 nsew signal output
rlabel metal2 s 96066 143200 96122 144000 6 wishbone_out[49]
port 530 nsew signal output
rlabel metal2 s 58622 143200 58678 144000 6 wishbone_out[4]
port 531 nsew signal output
rlabel metal2 s 96894 143200 96950 144000 6 wishbone_out[50]
port 532 nsew signal output
rlabel metal2 s 97722 143200 97778 144000 6 wishbone_out[51]
port 533 nsew signal output
rlabel metal2 s 98550 143200 98606 144000 6 wishbone_out[52]
port 534 nsew signal output
rlabel metal2 s 99378 143200 99434 144000 6 wishbone_out[53]
port 535 nsew signal output
rlabel metal2 s 100206 143200 100262 144000 6 wishbone_out[54]
port 536 nsew signal output
rlabel metal2 s 101034 143200 101090 144000 6 wishbone_out[55]
port 537 nsew signal output
rlabel metal2 s 101862 143200 101918 144000 6 wishbone_out[56]
port 538 nsew signal output
rlabel metal2 s 102690 143200 102746 144000 6 wishbone_out[57]
port 539 nsew signal output
rlabel metal2 s 103518 143200 103574 144000 6 wishbone_out[58]
port 540 nsew signal output
rlabel metal2 s 104346 143200 104402 144000 6 wishbone_out[59]
port 541 nsew signal output
rlabel metal2 s 59450 143200 59506 144000 6 wishbone_out[5]
port 542 nsew signal output
rlabel metal2 s 105174 143200 105230 144000 6 wishbone_out[60]
port 543 nsew signal output
rlabel metal2 s 106002 143200 106058 144000 6 wishbone_out[61]
port 544 nsew signal output
rlabel metal2 s 106830 143200 106886 144000 6 wishbone_out[62]
port 545 nsew signal output
rlabel metal2 s 107658 143200 107714 144000 6 wishbone_out[63]
port 546 nsew signal output
rlabel metal2 s 108578 143200 108634 144000 6 wishbone_out[64]
port 547 nsew signal output
rlabel metal2 s 109406 143200 109462 144000 6 wishbone_out[65]
port 548 nsew signal output
rlabel metal2 s 110234 143200 110290 144000 6 wishbone_out[66]
port 549 nsew signal output
rlabel metal2 s 111062 143200 111118 144000 6 wishbone_out[67]
port 550 nsew signal output
rlabel metal2 s 111890 143200 111946 144000 6 wishbone_out[68]
port 551 nsew signal output
rlabel metal2 s 112718 143200 112774 144000 6 wishbone_out[69]
port 552 nsew signal output
rlabel metal2 s 60278 143200 60334 144000 6 wishbone_out[6]
port 553 nsew signal output
rlabel metal2 s 113546 143200 113602 144000 6 wishbone_out[70]
port 554 nsew signal output
rlabel metal2 s 114374 143200 114430 144000 6 wishbone_out[71]
port 555 nsew signal output
rlabel metal2 s 115202 143200 115258 144000 6 wishbone_out[72]
port 556 nsew signal output
rlabel metal2 s 116030 143200 116086 144000 6 wishbone_out[73]
port 557 nsew signal output
rlabel metal2 s 116858 143200 116914 144000 6 wishbone_out[74]
port 558 nsew signal output
rlabel metal2 s 117686 143200 117742 144000 6 wishbone_out[75]
port 559 nsew signal output
rlabel metal2 s 118514 143200 118570 144000 6 wishbone_out[76]
port 560 nsew signal output
rlabel metal2 s 119342 143200 119398 144000 6 wishbone_out[77]
port 561 nsew signal output
rlabel metal2 s 120170 143200 120226 144000 6 wishbone_out[78]
port 562 nsew signal output
rlabel metal2 s 120998 143200 121054 144000 6 wishbone_out[79]
port 563 nsew signal output
rlabel metal2 s 61106 143200 61162 144000 6 wishbone_out[7]
port 564 nsew signal output
rlabel metal2 s 121826 143200 121882 144000 6 wishbone_out[80]
port 565 nsew signal output
rlabel metal2 s 122654 143200 122710 144000 6 wishbone_out[81]
port 566 nsew signal output
rlabel metal2 s 123482 143200 123538 144000 6 wishbone_out[82]
port 567 nsew signal output
rlabel metal2 s 124310 143200 124366 144000 6 wishbone_out[83]
port 568 nsew signal output
rlabel metal2 s 125138 143200 125194 144000 6 wishbone_out[84]
port 569 nsew signal output
rlabel metal2 s 125966 143200 126022 144000 6 wishbone_out[85]
port 570 nsew signal output
rlabel metal2 s 126886 143200 126942 144000 6 wishbone_out[86]
port 571 nsew signal output
rlabel metal2 s 127714 143200 127770 144000 6 wishbone_out[87]
port 572 nsew signal output
rlabel metal2 s 128542 143200 128598 144000 6 wishbone_out[88]
port 573 nsew signal output
rlabel metal2 s 129370 143200 129426 144000 6 wishbone_out[89]
port 574 nsew signal output
rlabel metal2 s 61934 143200 61990 144000 6 wishbone_out[8]
port 575 nsew signal output
rlabel metal2 s 130198 143200 130254 144000 6 wishbone_out[90]
port 576 nsew signal output
rlabel metal2 s 131026 143200 131082 144000 6 wishbone_out[91]
port 577 nsew signal output
rlabel metal2 s 131854 143200 131910 144000 6 wishbone_out[92]
port 578 nsew signal output
rlabel metal2 s 132682 143200 132738 144000 6 wishbone_out[93]
port 579 nsew signal output
rlabel metal2 s 133510 143200 133566 144000 6 wishbone_out[94]
port 580 nsew signal output
rlabel metal2 s 134338 143200 134394 144000 6 wishbone_out[95]
port 581 nsew signal output
rlabel metal2 s 135166 143200 135222 144000 6 wishbone_out[96]
port 582 nsew signal output
rlabel metal2 s 135994 143200 136050 144000 6 wishbone_out[97]
port 583 nsew signal output
rlabel metal2 s 136822 143200 136878 144000 6 wishbone_out[98]
port 584 nsew signal output
rlabel metal2 s 137650 143200 137706 144000 6 wishbone_out[99]
port 585 nsew signal output
rlabel metal2 s 62762 143200 62818 144000 6 wishbone_out[9]
port 586 nsew signal output
rlabel metal4 s 127088 2128 127408 141488 6 vccd1
port 587 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 141488 6 vccd1
port 588 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 141488 6 vccd1
port 589 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 141488 6 vccd1
port 590 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 141488 6 vccd1
port 591 nsew power bidirectional
rlabel metal4 s 111728 2128 112048 141488 6 vssd1
port 592 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 141488 6 vssd1
port 593 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 141488 6 vssd1
port 594 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 141488 6 vssd1
port 595 nsew ground bidirectional
rlabel metal4 s 127748 2176 128068 141440 6 vccd2
port 596 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 141440 6 vccd2
port 597 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 141440 6 vccd2
port 598 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 141440 6 vccd2
port 599 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 141440 6 vccd2
port 600 nsew power bidirectional
rlabel metal4 s 112388 2176 112708 141440 6 vssd2
port 601 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 141440 6 vssd2
port 602 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 141440 6 vssd2
port 603 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 141440 6 vssd2
port 604 nsew ground bidirectional
rlabel metal4 s 128408 2176 128728 141440 6 vdda1
port 605 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 141440 6 vdda1
port 606 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 141440 6 vdda1
port 607 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 141440 6 vdda1
port 608 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 141440 6 vdda1
port 609 nsew power bidirectional
rlabel metal4 s 113048 2176 113368 141440 6 vssa1
port 610 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 141440 6 vssa1
port 611 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 141440 6 vssa1
port 612 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 141440 6 vssa1
port 613 nsew ground bidirectional
rlabel metal4 s 129068 2176 129388 141440 6 vdda2
port 614 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 141440 6 vdda2
port 615 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 141440 6 vdda2
port 616 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 141440 6 vdda2
port 617 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 141440 6 vdda2
port 618 nsew power bidirectional
rlabel metal4 s 113708 2176 114028 141440 6 vssa2
port 619 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 141440 6 vssa2
port 620 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 141440 6 vssa2
port 621 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 141440 6 vssa2
port 622 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 143598 144000
string LEFview TRUE
<< end >>
