magic
tech sky130A
magscale 1 2
timestamp 1610960623
<< obsli1 >>
rect 866 2159 198821 197931
<< obsm1 >>
rect 144 348 199388 199980
<< metal2 >>
rect 148 199200 204 200000
rect 884 199200 940 200000
rect 1620 199200 1676 200000
rect 2448 199200 2504 200000
rect 3184 199200 3240 200000
rect 3920 199200 3976 200000
rect 4748 199200 4804 200000
rect 5484 199200 5540 200000
rect 6312 199200 6368 200000
rect 7048 199200 7104 200000
rect 7784 199200 7840 200000
rect 8612 199200 8668 200000
rect 9348 199200 9404 200000
rect 10176 199200 10232 200000
rect 10912 199200 10968 200000
rect 11648 199200 11704 200000
rect 12476 199200 12532 200000
rect 13212 199200 13268 200000
rect 14040 199200 14096 200000
rect 14776 199200 14832 200000
rect 15512 199200 15568 200000
rect 16340 199200 16396 200000
rect 17076 199200 17132 200000
rect 17904 199200 17960 200000
rect 18640 199200 18696 200000
rect 19376 199200 19432 200000
rect 20204 199200 20260 200000
rect 20940 199200 20996 200000
rect 21768 199200 21824 200000
rect 22504 199200 22560 200000
rect 23240 199200 23296 200000
rect 24068 199200 24124 200000
rect 24804 199200 24860 200000
rect 25540 199200 25596 200000
rect 26368 199200 26424 200000
rect 27104 199200 27160 200000
rect 27932 199200 27988 200000
rect 28668 199200 28724 200000
rect 29404 199200 29460 200000
rect 30232 199200 30288 200000
rect 30968 199200 31024 200000
rect 31796 199200 31852 200000
rect 32532 199200 32588 200000
rect 33268 199200 33324 200000
rect 34096 199200 34152 200000
rect 34832 199200 34888 200000
rect 35660 199200 35716 200000
rect 36396 199200 36452 200000
rect 37132 199200 37188 200000
rect 37960 199200 38016 200000
rect 38696 199200 38752 200000
rect 39524 199200 39580 200000
rect 40260 199200 40316 200000
rect 40996 199200 41052 200000
rect 41824 199200 41880 200000
rect 42560 199200 42616 200000
rect 43388 199200 43444 200000
rect 44124 199200 44180 200000
rect 44860 199200 44916 200000
rect 45688 199200 45744 200000
rect 46424 199200 46480 200000
rect 47252 199200 47308 200000
rect 47988 199200 48044 200000
rect 48724 199200 48780 200000
rect 49552 199200 49608 200000
rect 50288 199200 50344 200000
rect 51024 199200 51080 200000
rect 51852 199200 51908 200000
rect 52588 199200 52644 200000
rect 53416 199200 53472 200000
rect 54152 199200 54208 200000
rect 54888 199200 54944 200000
rect 55716 199200 55772 200000
rect 56452 199200 56508 200000
rect 57280 199200 57336 200000
rect 58016 199200 58072 200000
rect 58752 199200 58808 200000
rect 59580 199200 59636 200000
rect 60316 199200 60372 200000
rect 61144 199200 61200 200000
rect 61880 199200 61936 200000
rect 62616 199200 62672 200000
rect 63444 199200 63500 200000
rect 64180 199200 64236 200000
rect 65008 199200 65064 200000
rect 65744 199200 65800 200000
rect 66480 199200 66536 200000
rect 67308 199200 67364 200000
rect 68044 199200 68100 200000
rect 68872 199200 68928 200000
rect 69608 199200 69664 200000
rect 70344 199200 70400 200000
rect 71172 199200 71228 200000
rect 71908 199200 71964 200000
rect 72736 199200 72792 200000
rect 73472 199200 73528 200000
rect 74208 199200 74264 200000
rect 75036 199200 75092 200000
rect 75772 199200 75828 200000
rect 76508 199200 76564 200000
rect 77336 199200 77392 200000
rect 78072 199200 78128 200000
rect 78900 199200 78956 200000
rect 79636 199200 79692 200000
rect 80372 199200 80428 200000
rect 81200 199200 81256 200000
rect 81936 199200 81992 200000
rect 82764 199200 82820 200000
rect 83500 199200 83556 200000
rect 84236 199200 84292 200000
rect 85064 199200 85120 200000
rect 85800 199200 85856 200000
rect 86628 199200 86684 200000
rect 87364 199200 87420 200000
rect 88100 199200 88156 200000
rect 88928 199200 88984 200000
rect 89664 199200 89720 200000
rect 90492 199200 90548 200000
rect 91228 199200 91284 200000
rect 91964 199200 92020 200000
rect 92792 199200 92848 200000
rect 93528 199200 93584 200000
rect 94356 199200 94412 200000
rect 95092 199200 95148 200000
rect 95828 199200 95884 200000
rect 96656 199200 96712 200000
rect 97392 199200 97448 200000
rect 98220 199200 98276 200000
rect 98956 199200 99012 200000
rect 99692 199200 99748 200000
rect 100520 199200 100576 200000
rect 101256 199200 101312 200000
rect 101992 199200 102048 200000
rect 102820 199200 102876 200000
rect 103556 199200 103612 200000
rect 104384 199200 104440 200000
rect 105120 199200 105176 200000
rect 105856 199200 105912 200000
rect 106684 199200 106740 200000
rect 107420 199200 107476 200000
rect 108248 199200 108304 200000
rect 108984 199200 109040 200000
rect 109720 199200 109776 200000
rect 110548 199200 110604 200000
rect 111284 199200 111340 200000
rect 112112 199200 112168 200000
rect 112848 199200 112904 200000
rect 113584 199200 113640 200000
rect 114412 199200 114468 200000
rect 115148 199200 115204 200000
rect 115976 199200 116032 200000
rect 116712 199200 116768 200000
rect 117448 199200 117504 200000
rect 118276 199200 118332 200000
rect 119012 199200 119068 200000
rect 119840 199200 119896 200000
rect 120576 199200 120632 200000
rect 121312 199200 121368 200000
rect 122140 199200 122196 200000
rect 122876 199200 122932 200000
rect 123704 199200 123760 200000
rect 124440 199200 124496 200000
rect 125176 199200 125232 200000
rect 126004 199200 126060 200000
rect 126740 199200 126796 200000
rect 127476 199200 127532 200000
rect 128304 199200 128360 200000
rect 129040 199200 129096 200000
rect 129868 199200 129924 200000
rect 130604 199200 130660 200000
rect 131340 199200 131396 200000
rect 132168 199200 132224 200000
rect 132904 199200 132960 200000
rect 133732 199200 133788 200000
rect 134468 199200 134524 200000
rect 135204 199200 135260 200000
rect 136032 199200 136088 200000
rect 136768 199200 136824 200000
rect 137596 199200 137652 200000
rect 138332 199200 138388 200000
rect 139068 199200 139124 200000
rect 139896 199200 139952 200000
rect 140632 199200 140688 200000
rect 141460 199200 141516 200000
rect 142196 199200 142252 200000
rect 142932 199200 142988 200000
rect 143760 199200 143816 200000
rect 144496 199200 144552 200000
rect 145324 199200 145380 200000
rect 146060 199200 146116 200000
rect 146796 199200 146852 200000
rect 147624 199200 147680 200000
rect 148360 199200 148416 200000
rect 149188 199200 149244 200000
rect 149924 199200 149980 200000
rect 150660 199200 150716 200000
rect 151488 199200 151544 200000
rect 152224 199200 152280 200000
rect 152960 199200 153016 200000
rect 153788 199200 153844 200000
rect 154524 199200 154580 200000
rect 155352 199200 155408 200000
rect 156088 199200 156144 200000
rect 156824 199200 156880 200000
rect 157652 199200 157708 200000
rect 158388 199200 158444 200000
rect 159216 199200 159272 200000
rect 159952 199200 160008 200000
rect 160688 199200 160744 200000
rect 161516 199200 161572 200000
rect 162252 199200 162308 200000
rect 163080 199200 163136 200000
rect 163816 199200 163872 200000
rect 164552 199200 164608 200000
rect 165380 199200 165436 200000
rect 166116 199200 166172 200000
rect 166944 199200 167000 200000
rect 167680 199200 167736 200000
rect 168416 199200 168472 200000
rect 169244 199200 169300 200000
rect 169980 199200 170036 200000
rect 170808 199200 170864 200000
rect 171544 199200 171600 200000
rect 172280 199200 172336 200000
rect 173108 199200 173164 200000
rect 173844 199200 173900 200000
rect 174672 199200 174728 200000
rect 175408 199200 175464 200000
rect 176144 199200 176200 200000
rect 176972 199200 177028 200000
rect 177708 199200 177764 200000
rect 178444 199200 178500 200000
rect 179272 199200 179328 200000
rect 180008 199200 180064 200000
rect 180836 199200 180892 200000
rect 181572 199200 181628 200000
rect 182308 199200 182364 200000
rect 183136 199200 183192 200000
rect 183872 199200 183928 200000
rect 184700 199200 184756 200000
rect 185436 199200 185492 200000
rect 186172 199200 186228 200000
rect 187000 199200 187056 200000
rect 187736 199200 187792 200000
rect 188564 199200 188620 200000
rect 189300 199200 189356 200000
rect 190036 199200 190092 200000
rect 190864 199200 190920 200000
rect 191600 199200 191656 200000
rect 192428 199200 192484 200000
rect 193164 199200 193220 200000
rect 193900 199200 193956 200000
rect 194728 199200 194784 200000
rect 195464 199200 195520 200000
rect 196292 199200 196348 200000
rect 197028 199200 197084 200000
rect 197764 199200 197820 200000
rect 198592 199200 198648 200000
rect 199328 199200 199384 200000
rect 99784 0 99840 800
<< obsm2 >>
rect 56 199144 92 200025
rect 260 199144 828 200025
rect 996 199144 1564 200025
rect 1732 199144 2392 200025
rect 2560 199144 3128 200025
rect 3296 199144 3864 200025
rect 4032 199144 4692 200025
rect 4860 199144 5428 200025
rect 5596 199144 6256 200025
rect 6424 199144 6992 200025
rect 7160 199144 7728 200025
rect 7896 199144 8556 200025
rect 8724 199144 9292 200025
rect 9460 199144 10120 200025
rect 10288 199144 10856 200025
rect 11024 199144 11592 200025
rect 11760 199144 12420 200025
rect 12588 199144 13156 200025
rect 13324 199144 13984 200025
rect 14152 199144 14720 200025
rect 14888 199144 15456 200025
rect 15624 199144 16284 200025
rect 16452 199144 17020 200025
rect 17188 199144 17848 200025
rect 18016 199144 18584 200025
rect 18752 199144 19320 200025
rect 19488 199144 20148 200025
rect 20316 199144 20884 200025
rect 21052 199144 21712 200025
rect 21880 199144 22448 200025
rect 22616 199144 23184 200025
rect 23352 199144 24012 200025
rect 24180 199144 24748 200025
rect 24916 199144 25484 200025
rect 25652 199144 26312 200025
rect 26480 199144 27048 200025
rect 27216 199144 27876 200025
rect 28044 199144 28612 200025
rect 28780 199144 29348 200025
rect 29516 199144 30176 200025
rect 30344 199144 30912 200025
rect 31080 199144 31740 200025
rect 31908 199144 32476 200025
rect 32644 199144 33212 200025
rect 33380 199144 34040 200025
rect 34208 199144 34776 200025
rect 34944 199144 35604 200025
rect 35772 199144 36340 200025
rect 36508 199144 37076 200025
rect 37244 199144 37904 200025
rect 38072 199144 38640 200025
rect 38808 199144 39468 200025
rect 39636 199144 40204 200025
rect 40372 199144 40940 200025
rect 41108 199144 41768 200025
rect 41936 199144 42504 200025
rect 42672 199144 43332 200025
rect 43500 199144 44068 200025
rect 44236 199144 44804 200025
rect 44972 199144 45632 200025
rect 45800 199144 46368 200025
rect 46536 199144 47196 200025
rect 47364 199144 47932 200025
rect 48100 199144 48668 200025
rect 48836 199144 49496 200025
rect 49664 199144 50232 200025
rect 50400 199144 50968 200025
rect 51136 199144 51796 200025
rect 51964 199144 52532 200025
rect 52700 199144 53360 200025
rect 53528 199144 54096 200025
rect 54264 199144 54832 200025
rect 55000 199144 55660 200025
rect 55828 199144 56396 200025
rect 56564 199144 57224 200025
rect 57392 199144 57960 200025
rect 58128 199144 58696 200025
rect 58864 199144 59524 200025
rect 59692 199144 60260 200025
rect 60428 199144 61088 200025
rect 61256 199144 61824 200025
rect 61992 199144 62560 200025
rect 62728 199144 63388 200025
rect 63556 199144 64124 200025
rect 64292 199144 64952 200025
rect 65120 199144 65688 200025
rect 65856 199144 66424 200025
rect 66592 199144 67252 200025
rect 67420 199144 67988 200025
rect 68156 199144 68816 200025
rect 68984 199144 69552 200025
rect 69720 199144 70288 200025
rect 70456 199144 71116 200025
rect 71284 199144 71852 200025
rect 72020 199144 72680 200025
rect 72848 199144 73416 200025
rect 73584 199144 74152 200025
rect 74320 199144 74980 200025
rect 75148 199144 75716 200025
rect 75884 199144 76452 200025
rect 76620 199144 77280 200025
rect 77448 199144 78016 200025
rect 78184 199144 78844 200025
rect 79012 199144 79580 200025
rect 79748 199144 80316 200025
rect 80484 199144 81144 200025
rect 81312 199144 81880 200025
rect 82048 199144 82708 200025
rect 82876 199144 83444 200025
rect 83612 199144 84180 200025
rect 84348 199144 85008 200025
rect 85176 199144 85744 200025
rect 85912 199144 86572 200025
rect 86740 199144 87308 200025
rect 87476 199144 88044 200025
rect 88212 199144 88872 200025
rect 89040 199144 89608 200025
rect 89776 199144 90436 200025
rect 90604 199144 91172 200025
rect 91340 199144 91908 200025
rect 92076 199144 92736 200025
rect 92904 199144 93472 200025
rect 93640 199144 94300 200025
rect 94468 199144 95036 200025
rect 95204 199144 95772 200025
rect 95940 199144 96600 200025
rect 96768 199144 97336 200025
rect 97504 199144 98164 200025
rect 98332 199144 98900 200025
rect 99068 199144 99636 200025
rect 99804 199144 100464 200025
rect 100632 199144 101200 200025
rect 101368 199144 101936 200025
rect 102104 199144 102764 200025
rect 102932 199144 103500 200025
rect 103668 199144 104328 200025
rect 104496 199144 105064 200025
rect 105232 199144 105800 200025
rect 105968 199144 106628 200025
rect 106796 199144 107364 200025
rect 107532 199144 108192 200025
rect 108360 199144 108928 200025
rect 109096 199144 109664 200025
rect 109832 199144 110492 200025
rect 110660 199144 111228 200025
rect 111396 199144 112056 200025
rect 112224 199144 112792 200025
rect 112960 199144 113528 200025
rect 113696 199144 114356 200025
rect 114524 199144 115092 200025
rect 115260 199144 115920 200025
rect 116088 199144 116656 200025
rect 116824 199144 117392 200025
rect 117560 199144 118220 200025
rect 118388 199144 118956 200025
rect 119124 199144 119784 200025
rect 119952 199144 120520 200025
rect 120688 199144 121256 200025
rect 121424 199144 122084 200025
rect 122252 199144 122820 200025
rect 122988 199144 123648 200025
rect 123816 199144 124384 200025
rect 124552 199144 125120 200025
rect 125288 199144 125948 200025
rect 126116 199144 126684 200025
rect 126852 199144 127420 200025
rect 127588 199144 128248 200025
rect 128416 199144 128984 200025
rect 129152 199144 129812 200025
rect 129980 199144 130548 200025
rect 130716 199144 131284 200025
rect 131452 199144 132112 200025
rect 132280 199144 132848 200025
rect 133016 199144 133676 200025
rect 133844 199144 134412 200025
rect 134580 199144 135148 200025
rect 135316 199144 135976 200025
rect 136144 199144 136712 200025
rect 136880 199144 137540 200025
rect 137708 199144 138276 200025
rect 138444 199144 139012 200025
rect 139180 199144 139840 200025
rect 140008 199144 140576 200025
rect 140744 199144 141404 200025
rect 141572 199144 142140 200025
rect 142308 199144 142876 200025
rect 143044 199144 143704 200025
rect 143872 199144 144440 200025
rect 144608 199144 145268 200025
rect 145436 199144 146004 200025
rect 146172 199144 146740 200025
rect 146908 199144 147568 200025
rect 147736 199144 148304 200025
rect 148472 199144 149132 200025
rect 149300 199144 149868 200025
rect 150036 199144 150604 200025
rect 150772 199144 151432 200025
rect 151600 199144 152168 200025
rect 152336 199144 152904 200025
rect 153072 199144 153732 200025
rect 153900 199144 154468 200025
rect 154636 199144 155296 200025
rect 155464 199144 156032 200025
rect 156200 199144 156768 200025
rect 156936 199144 157596 200025
rect 157764 199144 158332 200025
rect 158500 199144 159160 200025
rect 159328 199144 159896 200025
rect 160064 199144 160632 200025
rect 160800 199144 161460 200025
rect 161628 199144 162196 200025
rect 162364 199144 163024 200025
rect 163192 199144 163760 200025
rect 163928 199144 164496 200025
rect 164664 199144 165324 200025
rect 165492 199144 166060 200025
rect 166228 199144 166888 200025
rect 167056 199144 167624 200025
rect 167792 199144 168360 200025
rect 168528 199144 169188 200025
rect 169356 199144 169924 200025
rect 170092 199144 170752 200025
rect 170920 199144 171488 200025
rect 171656 199144 172224 200025
rect 172392 199144 173052 200025
rect 173220 199144 173788 200025
rect 173956 199144 174616 200025
rect 174784 199144 175352 200025
rect 175520 199144 176088 200025
rect 176256 199144 176916 200025
rect 177084 199144 177652 200025
rect 177820 199144 178388 200025
rect 178556 199144 179216 200025
rect 179384 199144 179952 200025
rect 180120 199144 180780 200025
rect 180948 199144 181516 200025
rect 181684 199144 182252 200025
rect 182420 199144 183080 200025
rect 183248 199144 183816 200025
rect 183984 199144 184644 200025
rect 184812 199144 185380 200025
rect 185548 199144 186116 200025
rect 186284 199144 186944 200025
rect 187112 199144 187680 200025
rect 187848 199144 188508 200025
rect 188676 199144 189244 200025
rect 189412 199144 189980 200025
rect 190148 199144 190808 200025
rect 190976 199144 191544 200025
rect 191712 199144 192372 200025
rect 192540 199144 193108 200025
rect 193276 199144 193844 200025
rect 194012 199144 194672 200025
rect 194840 199144 195408 200025
rect 195576 199144 196236 200025
rect 196404 199144 196972 200025
rect 197140 199144 197708 200025
rect 197876 199144 198536 200025
rect 198704 199144 199272 200025
rect 56 856 199382 199144
rect 56 342 99728 856
rect 99896 342 199382 856
<< metal3 >>
rect 198962 199112 199762 199232
rect 198962 197616 199762 197736
rect 198962 196120 199762 196240
rect 198962 194488 199762 194608
rect 198962 192992 199762 193112
rect 198962 191496 199762 191616
rect 198962 189864 199762 189984
rect 198962 188368 199762 188488
rect 198962 186872 199762 186992
rect 198962 185240 199762 185360
rect 198962 183744 199762 183864
rect 198962 182248 199762 182368
rect 198962 180616 199762 180736
rect 198962 179120 199762 179240
rect 198962 177624 199762 177744
rect 198962 175992 199762 176112
rect 198962 174496 199762 174616
rect 198962 173000 199762 173120
rect 198962 171504 199762 171624
rect 198962 169872 199762 169992
rect 198962 168376 199762 168496
rect 198962 166880 199762 167000
rect 198962 165248 199762 165368
rect 198962 163752 199762 163872
rect 198962 162256 199762 162376
rect 198962 160624 199762 160744
rect 198962 159128 199762 159248
rect 198962 157632 199762 157752
rect 198962 156000 199762 156120
rect 198962 154504 199762 154624
rect 198962 153008 199762 153128
rect 198962 151376 199762 151496
rect 198962 149880 199762 150000
rect 198962 148384 199762 148504
rect 198962 146752 199762 146872
rect 198962 145256 199762 145376
rect 198962 143760 199762 143880
rect 198962 142264 199762 142384
rect 198962 140632 199762 140752
rect 198962 139136 199762 139256
rect 198962 137640 199762 137760
rect 198962 136008 199762 136128
rect 198962 134512 199762 134632
rect 198962 133016 199762 133136
rect 198962 131384 199762 131504
rect 198962 129888 199762 130008
rect 198962 128392 199762 128512
rect 198962 126760 199762 126880
rect 198962 125264 199762 125384
rect 198962 123768 199762 123888
rect 198962 122136 199762 122256
rect 198962 120640 199762 120760
rect 198962 119144 199762 119264
rect 198962 117512 199762 117632
rect 198962 116016 199762 116136
rect 198962 114520 199762 114640
rect 198962 113024 199762 113144
rect 198962 111392 199762 111512
rect 198962 109896 199762 110016
rect 198962 108400 199762 108520
rect 198962 106768 199762 106888
rect 198962 105272 199762 105392
rect 198962 103776 199762 103896
rect 198962 102144 199762 102264
rect 198962 100648 199762 100768
rect 198962 99152 199762 99272
rect 198962 97520 199762 97640
rect 198962 96024 199762 96144
rect 198962 94528 199762 94648
rect 198962 92896 199762 93016
rect 198962 91400 199762 91520
rect 198962 89904 199762 90024
rect 198962 88272 199762 88392
rect 198962 86776 199762 86896
rect 198962 85280 199762 85400
rect 198962 83784 199762 83904
rect 198962 82152 199762 82272
rect 198962 80656 199762 80776
rect 198962 79160 199762 79280
rect 198962 77528 199762 77648
rect 198962 76032 199762 76152
rect 198962 74536 199762 74656
rect 198962 72904 199762 73024
rect 198962 71408 199762 71528
rect 198962 69912 199762 70032
rect 198962 68280 199762 68400
rect 198962 66784 199762 66904
rect 198962 65288 199762 65408
rect 198962 63656 199762 63776
rect 198962 62160 199762 62280
rect 198962 60664 199762 60784
rect 198962 59032 199762 59152
rect 198962 57536 199762 57656
rect 198962 56040 199762 56160
rect 198962 54544 199762 54664
rect 198962 52912 199762 53032
rect 198962 51416 199762 51536
rect 198962 49920 199762 50040
rect 198962 48288 199762 48408
rect 198962 46792 199762 46912
rect 198962 45296 199762 45416
rect 198962 43664 199762 43784
rect 198962 42168 199762 42288
rect 198962 40672 199762 40792
rect 198962 39040 199762 39160
rect 198962 37544 199762 37664
rect 198962 36048 199762 36168
rect 198962 34416 199762 34536
rect 198962 32920 199762 33040
rect 198962 31424 199762 31544
rect 198962 29792 199762 29912
rect 198962 28296 199762 28416
rect 198962 26800 199762 26920
rect 198962 25304 199762 25424
rect 198962 23672 199762 23792
rect 198962 22176 199762 22296
rect 198962 20680 199762 20800
rect 198962 19048 199762 19168
rect 198962 17552 199762 17672
rect 198962 16056 199762 16176
rect 198962 14424 199762 14544
rect 198962 12928 199762 13048
rect 198962 11432 199762 11552
rect 198962 9800 199762 9920
rect 198962 8304 199762 8424
rect 198962 6808 199762 6928
rect 198962 5176 199762 5296
rect 198962 3680 199762 3800
rect 198962 2184 199762 2304
rect 198962 688 199762 808
<< obsm3 >>
rect 0 199312 199021 200021
rect 0 199032 198882 199312
rect 0 197816 199021 199032
rect 0 197536 198882 197816
rect 0 196320 199021 197536
rect 0 196040 198882 196320
rect 0 194688 199021 196040
rect 0 194408 198882 194688
rect 0 193192 199021 194408
rect 0 192912 198882 193192
rect 0 191696 199021 192912
rect 0 191416 198882 191696
rect 0 190064 199021 191416
rect 0 189784 198882 190064
rect 0 188568 199021 189784
rect 0 188288 198882 188568
rect 0 187072 199021 188288
rect 0 186792 198882 187072
rect 0 185440 199021 186792
rect 0 185160 198882 185440
rect 0 183944 199021 185160
rect 0 183664 198882 183944
rect 0 182448 199021 183664
rect 0 182168 198882 182448
rect 0 180816 199021 182168
rect 0 180536 198882 180816
rect 0 179320 199021 180536
rect 0 179040 198882 179320
rect 0 177824 199021 179040
rect 0 177544 198882 177824
rect 0 176192 199021 177544
rect 0 175912 198882 176192
rect 0 174696 199021 175912
rect 0 174416 198882 174696
rect 0 173200 199021 174416
rect 0 172920 198882 173200
rect 0 171704 199021 172920
rect 0 171424 198882 171704
rect 0 170072 199021 171424
rect 0 169792 198882 170072
rect 0 168576 199021 169792
rect 0 168296 198882 168576
rect 0 167080 199021 168296
rect 0 166800 198882 167080
rect 0 165448 199021 166800
rect 0 165168 198882 165448
rect 0 163952 199021 165168
rect 0 163672 198882 163952
rect 0 162456 199021 163672
rect 0 162176 198882 162456
rect 0 160824 199021 162176
rect 0 160544 198882 160824
rect 0 159328 199021 160544
rect 0 159048 198882 159328
rect 0 157832 199021 159048
rect 0 157552 198882 157832
rect 0 156200 199021 157552
rect 0 155920 198882 156200
rect 0 154704 199021 155920
rect 0 154424 198882 154704
rect 0 153208 199021 154424
rect 0 152928 198882 153208
rect 0 151576 199021 152928
rect 0 151296 198882 151576
rect 0 150080 199021 151296
rect 0 149800 198882 150080
rect 0 148584 199021 149800
rect 0 148304 198882 148584
rect 0 146952 199021 148304
rect 0 146672 198882 146952
rect 0 145456 199021 146672
rect 0 145176 198882 145456
rect 0 143960 199021 145176
rect 0 143680 198882 143960
rect 0 142464 199021 143680
rect 0 142184 198882 142464
rect 0 140832 199021 142184
rect 0 140552 198882 140832
rect 0 139336 199021 140552
rect 0 139056 198882 139336
rect 0 137840 199021 139056
rect 0 137560 198882 137840
rect 0 136208 199021 137560
rect 0 135928 198882 136208
rect 0 134712 199021 135928
rect 0 134432 198882 134712
rect 0 133216 199021 134432
rect 0 132936 198882 133216
rect 0 131584 199021 132936
rect 0 131304 198882 131584
rect 0 130088 199021 131304
rect 0 129808 198882 130088
rect 0 128592 199021 129808
rect 0 128312 198882 128592
rect 0 126960 199021 128312
rect 0 126680 198882 126960
rect 0 125464 199021 126680
rect 0 125184 198882 125464
rect 0 123968 199021 125184
rect 0 123688 198882 123968
rect 0 122336 199021 123688
rect 0 122056 198882 122336
rect 0 120840 199021 122056
rect 0 120560 198882 120840
rect 0 119344 199021 120560
rect 0 119064 198882 119344
rect 0 117712 199021 119064
rect 0 117432 198882 117712
rect 0 116216 199021 117432
rect 0 115936 198882 116216
rect 0 114720 199021 115936
rect 0 114440 198882 114720
rect 0 113224 199021 114440
rect 0 112944 198882 113224
rect 0 111592 199021 112944
rect 0 111312 198882 111592
rect 0 110096 199021 111312
rect 0 109816 198882 110096
rect 0 108600 199021 109816
rect 0 108320 198882 108600
rect 0 106968 199021 108320
rect 0 106688 198882 106968
rect 0 105472 199021 106688
rect 0 105192 198882 105472
rect 0 103976 199021 105192
rect 0 103696 198882 103976
rect 0 102344 199021 103696
rect 0 102064 198882 102344
rect 0 100848 199021 102064
rect 0 100568 198882 100848
rect 0 99352 199021 100568
rect 0 99072 198882 99352
rect 0 97720 199021 99072
rect 0 97440 198882 97720
rect 0 96224 199021 97440
rect 0 95944 198882 96224
rect 0 94728 199021 95944
rect 0 94448 198882 94728
rect 0 93096 199021 94448
rect 0 92816 198882 93096
rect 0 91600 199021 92816
rect 0 91320 198882 91600
rect 0 90104 199021 91320
rect 0 89824 198882 90104
rect 0 88472 199021 89824
rect 0 88192 198882 88472
rect 0 86976 199021 88192
rect 0 86696 198882 86976
rect 0 85480 199021 86696
rect 0 85200 198882 85480
rect 0 83984 199021 85200
rect 0 83704 198882 83984
rect 0 82352 199021 83704
rect 0 82072 198882 82352
rect 0 80856 199021 82072
rect 0 80576 198882 80856
rect 0 79360 199021 80576
rect 0 79080 198882 79360
rect 0 77728 199021 79080
rect 0 77448 198882 77728
rect 0 76232 199021 77448
rect 0 75952 198882 76232
rect 0 74736 199021 75952
rect 0 74456 198882 74736
rect 0 73104 199021 74456
rect 0 72824 198882 73104
rect 0 71608 199021 72824
rect 0 71328 198882 71608
rect 0 70112 199021 71328
rect 0 69832 198882 70112
rect 0 68480 199021 69832
rect 0 68200 198882 68480
rect 0 66984 199021 68200
rect 0 66704 198882 66984
rect 0 65488 199021 66704
rect 0 65208 198882 65488
rect 0 63856 199021 65208
rect 0 63576 198882 63856
rect 0 62360 199021 63576
rect 0 62080 198882 62360
rect 0 60864 199021 62080
rect 0 60584 198882 60864
rect 0 59232 199021 60584
rect 0 58952 198882 59232
rect 0 57736 199021 58952
rect 0 57456 198882 57736
rect 0 56240 199021 57456
rect 0 55960 198882 56240
rect 0 54744 199021 55960
rect 0 54464 198882 54744
rect 0 53112 199021 54464
rect 0 52832 198882 53112
rect 0 51616 199021 52832
rect 0 51336 198882 51616
rect 0 50120 199021 51336
rect 0 49840 198882 50120
rect 0 48488 199021 49840
rect 0 48208 198882 48488
rect 0 46992 199021 48208
rect 0 46712 198882 46992
rect 0 45496 199021 46712
rect 0 45216 198882 45496
rect 0 43864 199021 45216
rect 0 43584 198882 43864
rect 0 42368 199021 43584
rect 0 42088 198882 42368
rect 0 40872 199021 42088
rect 0 40592 198882 40872
rect 0 39240 199021 40592
rect 0 38960 198882 39240
rect 0 37744 199021 38960
rect 0 37464 198882 37744
rect 0 36248 199021 37464
rect 0 35968 198882 36248
rect 0 34616 199021 35968
rect 0 34336 198882 34616
rect 0 33120 199021 34336
rect 0 32840 198882 33120
rect 0 31624 199021 32840
rect 0 31344 198882 31624
rect 0 29992 199021 31344
rect 0 29712 198882 29992
rect 0 28496 199021 29712
rect 0 28216 198882 28496
rect 0 27000 199021 28216
rect 0 26720 198882 27000
rect 0 25504 199021 26720
rect 0 25224 198882 25504
rect 0 23872 199021 25224
rect 0 23592 198882 23872
rect 0 22376 199021 23592
rect 0 22096 198882 22376
rect 0 20880 199021 22096
rect 0 20600 198882 20880
rect 0 19248 199021 20600
rect 0 18968 198882 19248
rect 0 17752 199021 18968
rect 0 17472 198882 17752
rect 0 16256 199021 17472
rect 0 15976 198882 16256
rect 0 14624 199021 15976
rect 0 14344 198882 14624
rect 0 13128 199021 14344
rect 0 12848 198882 13128
rect 0 11632 199021 12848
rect 0 11352 198882 11632
rect 0 10000 199021 11352
rect 0 9720 198882 10000
rect 0 8504 199021 9720
rect 0 8224 198882 8504
rect 0 7008 199021 8224
rect 0 6728 198882 7008
rect 0 5376 199021 6728
rect 0 5096 198882 5376
rect 0 3880 199021 5096
rect 0 3600 198882 3880
rect 0 2384 199021 3600
rect 0 2104 198882 2384
rect 0 888 199021 2104
rect 0 608 198882 888
rect 0 579 199021 608
<< metal4 >>
rect 3970 2128 4290 197520
rect 4630 2176 4950 197472
rect 5290 2176 5610 197472
rect 5950 2176 6270 197472
rect 19330 2128 19650 197520
rect 19990 2176 20310 197472
rect 20650 2176 20970 197472
rect 21310 2176 21630 197472
rect 34690 2128 35010 197520
rect 35350 2176 35670 197472
rect 36010 2176 36330 197472
rect 36670 2176 36990 197472
rect 50050 2128 50370 197520
rect 50710 2176 51030 197472
rect 51370 2176 51690 197472
rect 52030 2176 52350 197472
rect 65410 2128 65730 197520
rect 66070 2176 66390 197472
rect 66730 2176 67050 197472
rect 67390 2176 67710 197472
rect 80770 2128 81090 197520
rect 81430 2176 81750 197472
rect 82090 2176 82410 197472
rect 82750 2176 83070 197472
rect 96130 2128 96450 197520
rect 96790 2176 97110 197472
rect 97450 2176 97770 197472
rect 98110 2176 98430 197472
rect 111490 2128 111810 197520
rect 112150 2176 112470 197472
rect 112810 2176 113130 197472
rect 113470 2176 113790 197472
rect 126850 2128 127170 197520
rect 127510 2176 127830 197472
rect 128170 2176 128490 197472
rect 128830 2176 129150 197472
rect 142210 2128 142530 197520
rect 142870 2176 143190 197472
rect 143530 2176 143850 197472
rect 144190 2176 144510 197472
rect 157570 2128 157890 197520
rect 158230 2176 158550 197472
rect 158890 2176 159210 197472
rect 159550 2176 159870 197472
rect 172930 2128 173250 197520
rect 173590 2176 173910 197472
rect 174250 2176 174570 197472
rect 174910 2176 175230 197472
rect 188290 2128 188610 197520
rect 188950 2176 189270 197472
rect 189610 2176 189930 197472
rect 190270 2176 190590 197472
<< obsm4 >>
rect 5 197600 196951 197981
rect 5 2048 3890 197600
rect 4370 197552 19250 197600
rect 4370 2096 4550 197552
rect 5030 2096 5210 197552
rect 5690 2096 5870 197552
rect 6350 2096 19250 197552
rect 19730 197552 34610 197600
rect 4370 2048 19250 2096
rect 19730 2096 19910 197552
rect 20390 2096 20570 197552
rect 21050 2096 21230 197552
rect 21710 2096 34610 197552
rect 35090 197552 49970 197600
rect 19730 2048 34610 2096
rect 35090 2096 35270 197552
rect 35750 2096 35930 197552
rect 36410 2096 36590 197552
rect 37070 2096 49970 197552
rect 50450 197552 65330 197600
rect 35090 2048 49970 2096
rect 50450 2096 50630 197552
rect 51110 2096 51290 197552
rect 51770 2096 51950 197552
rect 52430 2096 65330 197552
rect 65810 197552 80690 197600
rect 50450 2048 65330 2096
rect 65810 2096 65990 197552
rect 66470 2096 66650 197552
rect 67130 2096 67310 197552
rect 67790 2096 80690 197552
rect 81170 197552 96050 197600
rect 65810 2048 80690 2096
rect 81170 2096 81350 197552
rect 81830 2096 82010 197552
rect 82490 2096 82670 197552
rect 83150 2096 96050 197552
rect 96530 197552 111410 197600
rect 81170 2048 96050 2096
rect 96530 2096 96710 197552
rect 97190 2096 97370 197552
rect 97850 2096 98030 197552
rect 98510 2096 111410 197552
rect 111890 197552 126770 197600
rect 96530 2048 111410 2096
rect 111890 2096 112070 197552
rect 112550 2096 112730 197552
rect 113210 2096 113390 197552
rect 113870 2096 126770 197552
rect 127250 197552 142130 197600
rect 111890 2048 126770 2096
rect 127250 2096 127430 197552
rect 127910 2096 128090 197552
rect 128570 2096 128750 197552
rect 129230 2096 142130 197552
rect 142610 197552 157490 197600
rect 127250 2048 142130 2096
rect 142610 2096 142790 197552
rect 143270 2096 143450 197552
rect 143930 2096 144110 197552
rect 144590 2096 157490 197552
rect 157970 197552 172850 197600
rect 142610 2048 157490 2096
rect 157970 2096 158150 197552
rect 158630 2096 158810 197552
rect 159290 2096 159470 197552
rect 159950 2096 172850 197552
rect 173330 197552 188210 197600
rect 157970 2048 172850 2096
rect 173330 2096 173510 197552
rect 173990 2096 174170 197552
rect 174650 2096 174830 197552
rect 175310 2096 188210 197552
rect 188690 197552 196951 197600
rect 173330 2048 188210 2096
rect 188690 2096 188870 197552
rect 189350 2096 189530 197552
rect 190010 2096 190190 197552
rect 190670 2096 196951 197552
rect 188690 2048 196951 2096
rect 5 579 196951 2048
<< labels >>
rlabel metal2 s 99784 0 99840 800 6 clk
port 1 nsew signal input
rlabel metal2 s 148 199200 204 200000 6 m_in[0]
port 2 nsew signal input
rlabel metal2 s 77336 199200 77392 200000 6 m_in[100]
port 3 nsew signal input
rlabel metal2 s 78072 199200 78128 200000 6 m_in[101]
port 4 nsew signal input
rlabel metal2 s 78900 199200 78956 200000 6 m_in[102]
port 5 nsew signal input
rlabel metal2 s 79636 199200 79692 200000 6 m_in[103]
port 6 nsew signal input
rlabel metal2 s 80372 199200 80428 200000 6 m_in[104]
port 7 nsew signal input
rlabel metal2 s 81200 199200 81256 200000 6 m_in[105]
port 8 nsew signal input
rlabel metal2 s 81936 199200 81992 200000 6 m_in[106]
port 9 nsew signal input
rlabel metal2 s 82764 199200 82820 200000 6 m_in[107]
port 10 nsew signal input
rlabel metal2 s 83500 199200 83556 200000 6 m_in[108]
port 11 nsew signal input
rlabel metal2 s 84236 199200 84292 200000 6 m_in[109]
port 12 nsew signal input
rlabel metal2 s 7784 199200 7840 200000 6 m_in[10]
port 13 nsew signal input
rlabel metal2 s 85064 199200 85120 200000 6 m_in[110]
port 14 nsew signal input
rlabel metal2 s 85800 199200 85856 200000 6 m_in[111]
port 15 nsew signal input
rlabel metal2 s 86628 199200 86684 200000 6 m_in[112]
port 16 nsew signal input
rlabel metal2 s 87364 199200 87420 200000 6 m_in[113]
port 17 nsew signal input
rlabel metal2 s 88100 199200 88156 200000 6 m_in[114]
port 18 nsew signal input
rlabel metal2 s 88928 199200 88984 200000 6 m_in[115]
port 19 nsew signal input
rlabel metal2 s 89664 199200 89720 200000 6 m_in[116]
port 20 nsew signal input
rlabel metal2 s 90492 199200 90548 200000 6 m_in[117]
port 21 nsew signal input
rlabel metal2 s 91228 199200 91284 200000 6 m_in[118]
port 22 nsew signal input
rlabel metal2 s 91964 199200 92020 200000 6 m_in[119]
port 23 nsew signal input
rlabel metal2 s 8612 199200 8668 200000 6 m_in[11]
port 24 nsew signal input
rlabel metal2 s 92792 199200 92848 200000 6 m_in[120]
port 25 nsew signal input
rlabel metal2 s 93528 199200 93584 200000 6 m_in[121]
port 26 nsew signal input
rlabel metal2 s 94356 199200 94412 200000 6 m_in[122]
port 27 nsew signal input
rlabel metal2 s 95092 199200 95148 200000 6 m_in[123]
port 28 nsew signal input
rlabel metal2 s 95828 199200 95884 200000 6 m_in[124]
port 29 nsew signal input
rlabel metal2 s 96656 199200 96712 200000 6 m_in[125]
port 30 nsew signal input
rlabel metal2 s 97392 199200 97448 200000 6 m_in[126]
port 31 nsew signal input
rlabel metal2 s 98220 199200 98276 200000 6 m_in[127]
port 32 nsew signal input
rlabel metal2 s 98956 199200 99012 200000 6 m_in[128]
port 33 nsew signal input
rlabel metal2 s 99692 199200 99748 200000 6 m_in[129]
port 34 nsew signal input
rlabel metal2 s 9348 199200 9404 200000 6 m_in[12]
port 35 nsew signal input
rlabel metal2 s 100520 199200 100576 200000 6 m_in[130]
port 36 nsew signal input
rlabel metal2 s 101256 199200 101312 200000 6 m_in[131]
port 37 nsew signal input
rlabel metal2 s 101992 199200 102048 200000 6 m_in[132]
port 38 nsew signal input
rlabel metal2 s 102820 199200 102876 200000 6 m_in[133]
port 39 nsew signal input
rlabel metal2 s 103556 199200 103612 200000 6 m_in[134]
port 40 nsew signal input
rlabel metal2 s 104384 199200 104440 200000 6 m_in[135]
port 41 nsew signal input
rlabel metal2 s 105120 199200 105176 200000 6 m_in[136]
port 42 nsew signal input
rlabel metal2 s 105856 199200 105912 200000 6 m_in[137]
port 43 nsew signal input
rlabel metal2 s 106684 199200 106740 200000 6 m_in[138]
port 44 nsew signal input
rlabel metal2 s 107420 199200 107476 200000 6 m_in[139]
port 45 nsew signal input
rlabel metal2 s 10176 199200 10232 200000 6 m_in[13]
port 46 nsew signal input
rlabel metal2 s 108248 199200 108304 200000 6 m_in[140]
port 47 nsew signal input
rlabel metal2 s 108984 199200 109040 200000 6 m_in[141]
port 48 nsew signal input
rlabel metal2 s 109720 199200 109776 200000 6 m_in[142]
port 49 nsew signal input
rlabel metal2 s 110548 199200 110604 200000 6 m_in[143]
port 50 nsew signal input
rlabel metal2 s 111284 199200 111340 200000 6 m_in[144]
port 51 nsew signal input
rlabel metal2 s 112112 199200 112168 200000 6 m_in[145]
port 52 nsew signal input
rlabel metal2 s 112848 199200 112904 200000 6 m_in[146]
port 53 nsew signal input
rlabel metal2 s 113584 199200 113640 200000 6 m_in[147]
port 54 nsew signal input
rlabel metal2 s 114412 199200 114468 200000 6 m_in[148]
port 55 nsew signal input
rlabel metal2 s 115148 199200 115204 200000 6 m_in[149]
port 56 nsew signal input
rlabel metal2 s 10912 199200 10968 200000 6 m_in[14]
port 57 nsew signal input
rlabel metal2 s 115976 199200 116032 200000 6 m_in[150]
port 58 nsew signal input
rlabel metal2 s 116712 199200 116768 200000 6 m_in[151]
port 59 nsew signal input
rlabel metal2 s 117448 199200 117504 200000 6 m_in[152]
port 60 nsew signal input
rlabel metal2 s 118276 199200 118332 200000 6 m_in[153]
port 61 nsew signal input
rlabel metal2 s 119012 199200 119068 200000 6 m_in[154]
port 62 nsew signal input
rlabel metal2 s 119840 199200 119896 200000 6 m_in[155]
port 63 nsew signal input
rlabel metal2 s 120576 199200 120632 200000 6 m_in[156]
port 64 nsew signal input
rlabel metal2 s 121312 199200 121368 200000 6 m_in[157]
port 65 nsew signal input
rlabel metal2 s 122140 199200 122196 200000 6 m_in[158]
port 66 nsew signal input
rlabel metal2 s 122876 199200 122932 200000 6 m_in[159]
port 67 nsew signal input
rlabel metal2 s 11648 199200 11704 200000 6 m_in[15]
port 68 nsew signal input
rlabel metal2 s 123704 199200 123760 200000 6 m_in[160]
port 69 nsew signal input
rlabel metal2 s 124440 199200 124496 200000 6 m_in[161]
port 70 nsew signal input
rlabel metal2 s 125176 199200 125232 200000 6 m_in[162]
port 71 nsew signal input
rlabel metal2 s 126004 199200 126060 200000 6 m_in[163]
port 72 nsew signal input
rlabel metal2 s 126740 199200 126796 200000 6 m_in[164]
port 73 nsew signal input
rlabel metal2 s 127476 199200 127532 200000 6 m_in[165]
port 74 nsew signal input
rlabel metal2 s 128304 199200 128360 200000 6 m_in[166]
port 75 nsew signal input
rlabel metal2 s 129040 199200 129096 200000 6 m_in[167]
port 76 nsew signal input
rlabel metal2 s 129868 199200 129924 200000 6 m_in[168]
port 77 nsew signal input
rlabel metal2 s 130604 199200 130660 200000 6 m_in[169]
port 78 nsew signal input
rlabel metal2 s 12476 199200 12532 200000 6 m_in[16]
port 79 nsew signal input
rlabel metal2 s 131340 199200 131396 200000 6 m_in[170]
port 80 nsew signal input
rlabel metal2 s 132168 199200 132224 200000 6 m_in[171]
port 81 nsew signal input
rlabel metal2 s 132904 199200 132960 200000 6 m_in[172]
port 82 nsew signal input
rlabel metal2 s 133732 199200 133788 200000 6 m_in[173]
port 83 nsew signal input
rlabel metal2 s 134468 199200 134524 200000 6 m_in[174]
port 84 nsew signal input
rlabel metal2 s 135204 199200 135260 200000 6 m_in[175]
port 85 nsew signal input
rlabel metal2 s 136032 199200 136088 200000 6 m_in[176]
port 86 nsew signal input
rlabel metal2 s 136768 199200 136824 200000 6 m_in[177]
port 87 nsew signal input
rlabel metal2 s 137596 199200 137652 200000 6 m_in[178]
port 88 nsew signal input
rlabel metal2 s 138332 199200 138388 200000 6 m_in[179]
port 89 nsew signal input
rlabel metal2 s 13212 199200 13268 200000 6 m_in[17]
port 90 nsew signal input
rlabel metal2 s 139068 199200 139124 200000 6 m_in[180]
port 91 nsew signal input
rlabel metal2 s 139896 199200 139952 200000 6 m_in[181]
port 92 nsew signal input
rlabel metal2 s 140632 199200 140688 200000 6 m_in[182]
port 93 nsew signal input
rlabel metal2 s 141460 199200 141516 200000 6 m_in[183]
port 94 nsew signal input
rlabel metal2 s 142196 199200 142252 200000 6 m_in[184]
port 95 nsew signal input
rlabel metal2 s 142932 199200 142988 200000 6 m_in[185]
port 96 nsew signal input
rlabel metal2 s 143760 199200 143816 200000 6 m_in[186]
port 97 nsew signal input
rlabel metal2 s 144496 199200 144552 200000 6 m_in[187]
port 98 nsew signal input
rlabel metal2 s 145324 199200 145380 200000 6 m_in[188]
port 99 nsew signal input
rlabel metal2 s 146060 199200 146116 200000 6 m_in[189]
port 100 nsew signal input
rlabel metal2 s 14040 199200 14096 200000 6 m_in[18]
port 101 nsew signal input
rlabel metal2 s 146796 199200 146852 200000 6 m_in[190]
port 102 nsew signal input
rlabel metal2 s 147624 199200 147680 200000 6 m_in[191]
port 103 nsew signal input
rlabel metal2 s 148360 199200 148416 200000 6 m_in[192]
port 104 nsew signal input
rlabel metal2 s 149188 199200 149244 200000 6 m_in[193]
port 105 nsew signal input
rlabel metal2 s 149924 199200 149980 200000 6 m_in[194]
port 106 nsew signal input
rlabel metal2 s 150660 199200 150716 200000 6 m_in[195]
port 107 nsew signal input
rlabel metal2 s 151488 199200 151544 200000 6 m_in[196]
port 108 nsew signal input
rlabel metal2 s 152224 199200 152280 200000 6 m_in[197]
port 109 nsew signal input
rlabel metal2 s 152960 199200 153016 200000 6 m_in[198]
port 110 nsew signal input
rlabel metal2 s 153788 199200 153844 200000 6 m_in[199]
port 111 nsew signal input
rlabel metal2 s 14776 199200 14832 200000 6 m_in[19]
port 112 nsew signal input
rlabel metal2 s 884 199200 940 200000 6 m_in[1]
port 113 nsew signal input
rlabel metal2 s 154524 199200 154580 200000 6 m_in[200]
port 114 nsew signal input
rlabel metal2 s 155352 199200 155408 200000 6 m_in[201]
port 115 nsew signal input
rlabel metal2 s 156088 199200 156144 200000 6 m_in[202]
port 116 nsew signal input
rlabel metal2 s 156824 199200 156880 200000 6 m_in[203]
port 117 nsew signal input
rlabel metal2 s 157652 199200 157708 200000 6 m_in[204]
port 118 nsew signal input
rlabel metal2 s 158388 199200 158444 200000 6 m_in[205]
port 119 nsew signal input
rlabel metal2 s 159216 199200 159272 200000 6 m_in[206]
port 120 nsew signal input
rlabel metal2 s 159952 199200 160008 200000 6 m_in[207]
port 121 nsew signal input
rlabel metal2 s 160688 199200 160744 200000 6 m_in[208]
port 122 nsew signal input
rlabel metal2 s 161516 199200 161572 200000 6 m_in[209]
port 123 nsew signal input
rlabel metal2 s 15512 199200 15568 200000 6 m_in[20]
port 124 nsew signal input
rlabel metal2 s 162252 199200 162308 200000 6 m_in[210]
port 125 nsew signal input
rlabel metal2 s 163080 199200 163136 200000 6 m_in[211]
port 126 nsew signal input
rlabel metal2 s 163816 199200 163872 200000 6 m_in[212]
port 127 nsew signal input
rlabel metal2 s 164552 199200 164608 200000 6 m_in[213]
port 128 nsew signal input
rlabel metal2 s 165380 199200 165436 200000 6 m_in[214]
port 129 nsew signal input
rlabel metal2 s 166116 199200 166172 200000 6 m_in[215]
port 130 nsew signal input
rlabel metal2 s 166944 199200 167000 200000 6 m_in[216]
port 131 nsew signal input
rlabel metal2 s 167680 199200 167736 200000 6 m_in[217]
port 132 nsew signal input
rlabel metal2 s 168416 199200 168472 200000 6 m_in[218]
port 133 nsew signal input
rlabel metal2 s 169244 199200 169300 200000 6 m_in[219]
port 134 nsew signal input
rlabel metal2 s 16340 199200 16396 200000 6 m_in[21]
port 135 nsew signal input
rlabel metal2 s 169980 199200 170036 200000 6 m_in[220]
port 136 nsew signal input
rlabel metal2 s 170808 199200 170864 200000 6 m_in[221]
port 137 nsew signal input
rlabel metal2 s 171544 199200 171600 200000 6 m_in[222]
port 138 nsew signal input
rlabel metal2 s 172280 199200 172336 200000 6 m_in[223]
port 139 nsew signal input
rlabel metal2 s 173108 199200 173164 200000 6 m_in[224]
port 140 nsew signal input
rlabel metal2 s 173844 199200 173900 200000 6 m_in[225]
port 141 nsew signal input
rlabel metal2 s 174672 199200 174728 200000 6 m_in[226]
port 142 nsew signal input
rlabel metal2 s 175408 199200 175464 200000 6 m_in[227]
port 143 nsew signal input
rlabel metal2 s 176144 199200 176200 200000 6 m_in[228]
port 144 nsew signal input
rlabel metal2 s 176972 199200 177028 200000 6 m_in[229]
port 145 nsew signal input
rlabel metal2 s 17076 199200 17132 200000 6 m_in[22]
port 146 nsew signal input
rlabel metal2 s 177708 199200 177764 200000 6 m_in[230]
port 147 nsew signal input
rlabel metal2 s 178444 199200 178500 200000 6 m_in[231]
port 148 nsew signal input
rlabel metal2 s 179272 199200 179328 200000 6 m_in[232]
port 149 nsew signal input
rlabel metal2 s 180008 199200 180064 200000 6 m_in[233]
port 150 nsew signal input
rlabel metal2 s 180836 199200 180892 200000 6 m_in[234]
port 151 nsew signal input
rlabel metal2 s 181572 199200 181628 200000 6 m_in[235]
port 152 nsew signal input
rlabel metal2 s 182308 199200 182364 200000 6 m_in[236]
port 153 nsew signal input
rlabel metal2 s 183136 199200 183192 200000 6 m_in[237]
port 154 nsew signal input
rlabel metal2 s 183872 199200 183928 200000 6 m_in[238]
port 155 nsew signal input
rlabel metal2 s 184700 199200 184756 200000 6 m_in[239]
port 156 nsew signal input
rlabel metal2 s 17904 199200 17960 200000 6 m_in[23]
port 157 nsew signal input
rlabel metal2 s 185436 199200 185492 200000 6 m_in[240]
port 158 nsew signal input
rlabel metal2 s 186172 199200 186228 200000 6 m_in[241]
port 159 nsew signal input
rlabel metal2 s 187000 199200 187056 200000 6 m_in[242]
port 160 nsew signal input
rlabel metal2 s 187736 199200 187792 200000 6 m_in[243]
port 161 nsew signal input
rlabel metal2 s 188564 199200 188620 200000 6 m_in[244]
port 162 nsew signal input
rlabel metal2 s 189300 199200 189356 200000 6 m_in[245]
port 163 nsew signal input
rlabel metal2 s 190036 199200 190092 200000 6 m_in[246]
port 164 nsew signal input
rlabel metal2 s 190864 199200 190920 200000 6 m_in[247]
port 165 nsew signal input
rlabel metal2 s 191600 199200 191656 200000 6 m_in[248]
port 166 nsew signal input
rlabel metal2 s 192428 199200 192484 200000 6 m_in[249]
port 167 nsew signal input
rlabel metal2 s 18640 199200 18696 200000 6 m_in[24]
port 168 nsew signal input
rlabel metal2 s 193164 199200 193220 200000 6 m_in[250]
port 169 nsew signal input
rlabel metal2 s 193900 199200 193956 200000 6 m_in[251]
port 170 nsew signal input
rlabel metal2 s 194728 199200 194784 200000 6 m_in[252]
port 171 nsew signal input
rlabel metal2 s 195464 199200 195520 200000 6 m_in[253]
port 172 nsew signal input
rlabel metal2 s 196292 199200 196348 200000 6 m_in[254]
port 173 nsew signal input
rlabel metal2 s 197028 199200 197084 200000 6 m_in[255]
port 174 nsew signal input
rlabel metal2 s 197764 199200 197820 200000 6 m_in[256]
port 175 nsew signal input
rlabel metal2 s 198592 199200 198648 200000 6 m_in[257]
port 176 nsew signal input
rlabel metal2 s 199328 199200 199384 200000 6 m_in[258]
port 177 nsew signal input
rlabel metal2 s 19376 199200 19432 200000 6 m_in[25]
port 178 nsew signal input
rlabel metal2 s 20204 199200 20260 200000 6 m_in[26]
port 179 nsew signal input
rlabel metal2 s 20940 199200 20996 200000 6 m_in[27]
port 180 nsew signal input
rlabel metal2 s 21768 199200 21824 200000 6 m_in[28]
port 181 nsew signal input
rlabel metal2 s 22504 199200 22560 200000 6 m_in[29]
port 182 nsew signal input
rlabel metal2 s 1620 199200 1676 200000 6 m_in[2]
port 183 nsew signal input
rlabel metal2 s 23240 199200 23296 200000 6 m_in[30]
port 184 nsew signal input
rlabel metal2 s 24068 199200 24124 200000 6 m_in[31]
port 185 nsew signal input
rlabel metal2 s 24804 199200 24860 200000 6 m_in[32]
port 186 nsew signal input
rlabel metal2 s 25540 199200 25596 200000 6 m_in[33]
port 187 nsew signal input
rlabel metal2 s 26368 199200 26424 200000 6 m_in[34]
port 188 nsew signal input
rlabel metal2 s 27104 199200 27160 200000 6 m_in[35]
port 189 nsew signal input
rlabel metal2 s 27932 199200 27988 200000 6 m_in[36]
port 190 nsew signal input
rlabel metal2 s 28668 199200 28724 200000 6 m_in[37]
port 191 nsew signal input
rlabel metal2 s 29404 199200 29460 200000 6 m_in[38]
port 192 nsew signal input
rlabel metal2 s 30232 199200 30288 200000 6 m_in[39]
port 193 nsew signal input
rlabel metal2 s 2448 199200 2504 200000 6 m_in[3]
port 194 nsew signal input
rlabel metal2 s 30968 199200 31024 200000 6 m_in[40]
port 195 nsew signal input
rlabel metal2 s 31796 199200 31852 200000 6 m_in[41]
port 196 nsew signal input
rlabel metal2 s 32532 199200 32588 200000 6 m_in[42]
port 197 nsew signal input
rlabel metal2 s 33268 199200 33324 200000 6 m_in[43]
port 198 nsew signal input
rlabel metal2 s 34096 199200 34152 200000 6 m_in[44]
port 199 nsew signal input
rlabel metal2 s 34832 199200 34888 200000 6 m_in[45]
port 200 nsew signal input
rlabel metal2 s 35660 199200 35716 200000 6 m_in[46]
port 201 nsew signal input
rlabel metal2 s 36396 199200 36452 200000 6 m_in[47]
port 202 nsew signal input
rlabel metal2 s 37132 199200 37188 200000 6 m_in[48]
port 203 nsew signal input
rlabel metal2 s 37960 199200 38016 200000 6 m_in[49]
port 204 nsew signal input
rlabel metal2 s 3184 199200 3240 200000 6 m_in[4]
port 205 nsew signal input
rlabel metal2 s 38696 199200 38752 200000 6 m_in[50]
port 206 nsew signal input
rlabel metal2 s 39524 199200 39580 200000 6 m_in[51]
port 207 nsew signal input
rlabel metal2 s 40260 199200 40316 200000 6 m_in[52]
port 208 nsew signal input
rlabel metal2 s 40996 199200 41052 200000 6 m_in[53]
port 209 nsew signal input
rlabel metal2 s 41824 199200 41880 200000 6 m_in[54]
port 210 nsew signal input
rlabel metal2 s 42560 199200 42616 200000 6 m_in[55]
port 211 nsew signal input
rlabel metal2 s 43388 199200 43444 200000 6 m_in[56]
port 212 nsew signal input
rlabel metal2 s 44124 199200 44180 200000 6 m_in[57]
port 213 nsew signal input
rlabel metal2 s 44860 199200 44916 200000 6 m_in[58]
port 214 nsew signal input
rlabel metal2 s 45688 199200 45744 200000 6 m_in[59]
port 215 nsew signal input
rlabel metal2 s 3920 199200 3976 200000 6 m_in[5]
port 216 nsew signal input
rlabel metal2 s 46424 199200 46480 200000 6 m_in[60]
port 217 nsew signal input
rlabel metal2 s 47252 199200 47308 200000 6 m_in[61]
port 218 nsew signal input
rlabel metal2 s 47988 199200 48044 200000 6 m_in[62]
port 219 nsew signal input
rlabel metal2 s 48724 199200 48780 200000 6 m_in[63]
port 220 nsew signal input
rlabel metal2 s 49552 199200 49608 200000 6 m_in[64]
port 221 nsew signal input
rlabel metal2 s 50288 199200 50344 200000 6 m_in[65]
port 222 nsew signal input
rlabel metal2 s 51024 199200 51080 200000 6 m_in[66]
port 223 nsew signal input
rlabel metal2 s 51852 199200 51908 200000 6 m_in[67]
port 224 nsew signal input
rlabel metal2 s 52588 199200 52644 200000 6 m_in[68]
port 225 nsew signal input
rlabel metal2 s 53416 199200 53472 200000 6 m_in[69]
port 226 nsew signal input
rlabel metal2 s 4748 199200 4804 200000 6 m_in[6]
port 227 nsew signal input
rlabel metal2 s 54152 199200 54208 200000 6 m_in[70]
port 228 nsew signal input
rlabel metal2 s 54888 199200 54944 200000 6 m_in[71]
port 229 nsew signal input
rlabel metal2 s 55716 199200 55772 200000 6 m_in[72]
port 230 nsew signal input
rlabel metal2 s 56452 199200 56508 200000 6 m_in[73]
port 231 nsew signal input
rlabel metal2 s 57280 199200 57336 200000 6 m_in[74]
port 232 nsew signal input
rlabel metal2 s 58016 199200 58072 200000 6 m_in[75]
port 233 nsew signal input
rlabel metal2 s 58752 199200 58808 200000 6 m_in[76]
port 234 nsew signal input
rlabel metal2 s 59580 199200 59636 200000 6 m_in[77]
port 235 nsew signal input
rlabel metal2 s 60316 199200 60372 200000 6 m_in[78]
port 236 nsew signal input
rlabel metal2 s 61144 199200 61200 200000 6 m_in[79]
port 237 nsew signal input
rlabel metal2 s 5484 199200 5540 200000 6 m_in[7]
port 238 nsew signal input
rlabel metal2 s 61880 199200 61936 200000 6 m_in[80]
port 239 nsew signal input
rlabel metal2 s 62616 199200 62672 200000 6 m_in[81]
port 240 nsew signal input
rlabel metal2 s 63444 199200 63500 200000 6 m_in[82]
port 241 nsew signal input
rlabel metal2 s 64180 199200 64236 200000 6 m_in[83]
port 242 nsew signal input
rlabel metal2 s 65008 199200 65064 200000 6 m_in[84]
port 243 nsew signal input
rlabel metal2 s 65744 199200 65800 200000 6 m_in[85]
port 244 nsew signal input
rlabel metal2 s 66480 199200 66536 200000 6 m_in[86]
port 245 nsew signal input
rlabel metal2 s 67308 199200 67364 200000 6 m_in[87]
port 246 nsew signal input
rlabel metal2 s 68044 199200 68100 200000 6 m_in[88]
port 247 nsew signal input
rlabel metal2 s 68872 199200 68928 200000 6 m_in[89]
port 248 nsew signal input
rlabel metal2 s 6312 199200 6368 200000 6 m_in[8]
port 249 nsew signal input
rlabel metal2 s 69608 199200 69664 200000 6 m_in[90]
port 250 nsew signal input
rlabel metal2 s 70344 199200 70400 200000 6 m_in[91]
port 251 nsew signal input
rlabel metal2 s 71172 199200 71228 200000 6 m_in[92]
port 252 nsew signal input
rlabel metal2 s 71908 199200 71964 200000 6 m_in[93]
port 253 nsew signal input
rlabel metal2 s 72736 199200 72792 200000 6 m_in[94]
port 254 nsew signal input
rlabel metal2 s 73472 199200 73528 200000 6 m_in[95]
port 255 nsew signal input
rlabel metal2 s 74208 199200 74264 200000 6 m_in[96]
port 256 nsew signal input
rlabel metal2 s 75036 199200 75092 200000 6 m_in[97]
port 257 nsew signal input
rlabel metal2 s 75772 199200 75828 200000 6 m_in[98]
port 258 nsew signal input
rlabel metal2 s 76508 199200 76564 200000 6 m_in[99]
port 259 nsew signal input
rlabel metal2 s 7048 199200 7104 200000 6 m_in[9]
port 260 nsew signal input
rlabel metal3 s 198962 688 199762 808 6 m_out[0]
port 261 nsew signal output
rlabel metal3 s 198962 154504 199762 154624 6 m_out[100]
port 262 nsew signal output
rlabel metal3 s 198962 156000 199762 156120 6 m_out[101]
port 263 nsew signal output
rlabel metal3 s 198962 157632 199762 157752 6 m_out[102]
port 264 nsew signal output
rlabel metal3 s 198962 159128 199762 159248 6 m_out[103]
port 265 nsew signal output
rlabel metal3 s 198962 160624 199762 160744 6 m_out[104]
port 266 nsew signal output
rlabel metal3 s 198962 162256 199762 162376 6 m_out[105]
port 267 nsew signal output
rlabel metal3 s 198962 163752 199762 163872 6 m_out[106]
port 268 nsew signal output
rlabel metal3 s 198962 165248 199762 165368 6 m_out[107]
port 269 nsew signal output
rlabel metal3 s 198962 166880 199762 167000 6 m_out[108]
port 270 nsew signal output
rlabel metal3 s 198962 168376 199762 168496 6 m_out[109]
port 271 nsew signal output
rlabel metal3 s 198962 16056 199762 16176 6 m_out[10]
port 272 nsew signal output
rlabel metal3 s 198962 169872 199762 169992 6 m_out[110]
port 273 nsew signal output
rlabel metal3 s 198962 171504 199762 171624 6 m_out[111]
port 274 nsew signal output
rlabel metal3 s 198962 173000 199762 173120 6 m_out[112]
port 275 nsew signal output
rlabel metal3 s 198962 174496 199762 174616 6 m_out[113]
port 276 nsew signal output
rlabel metal3 s 198962 175992 199762 176112 6 m_out[114]
port 277 nsew signal output
rlabel metal3 s 198962 177624 199762 177744 6 m_out[115]
port 278 nsew signal output
rlabel metal3 s 198962 179120 199762 179240 6 m_out[116]
port 279 nsew signal output
rlabel metal3 s 198962 180616 199762 180736 6 m_out[117]
port 280 nsew signal output
rlabel metal3 s 198962 182248 199762 182368 6 m_out[118]
port 281 nsew signal output
rlabel metal3 s 198962 183744 199762 183864 6 m_out[119]
port 282 nsew signal output
rlabel metal3 s 198962 17552 199762 17672 6 m_out[11]
port 283 nsew signal output
rlabel metal3 s 198962 185240 199762 185360 6 m_out[120]
port 284 nsew signal output
rlabel metal3 s 198962 186872 199762 186992 6 m_out[121]
port 285 nsew signal output
rlabel metal3 s 198962 188368 199762 188488 6 m_out[122]
port 286 nsew signal output
rlabel metal3 s 198962 189864 199762 189984 6 m_out[123]
port 287 nsew signal output
rlabel metal3 s 198962 191496 199762 191616 6 m_out[124]
port 288 nsew signal output
rlabel metal3 s 198962 192992 199762 193112 6 m_out[125]
port 289 nsew signal output
rlabel metal3 s 198962 194488 199762 194608 6 m_out[126]
port 290 nsew signal output
rlabel metal3 s 198962 196120 199762 196240 6 m_out[127]
port 291 nsew signal output
rlabel metal3 s 198962 197616 199762 197736 6 m_out[128]
port 292 nsew signal output
rlabel metal3 s 198962 199112 199762 199232 6 m_out[129]
port 293 nsew signal output
rlabel metal3 s 198962 19048 199762 19168 6 m_out[12]
port 294 nsew signal output
rlabel metal3 s 198962 20680 199762 20800 6 m_out[13]
port 295 nsew signal output
rlabel metal3 s 198962 22176 199762 22296 6 m_out[14]
port 296 nsew signal output
rlabel metal3 s 198962 23672 199762 23792 6 m_out[15]
port 297 nsew signal output
rlabel metal3 s 198962 25304 199762 25424 6 m_out[16]
port 298 nsew signal output
rlabel metal3 s 198962 26800 199762 26920 6 m_out[17]
port 299 nsew signal output
rlabel metal3 s 198962 28296 199762 28416 6 m_out[18]
port 300 nsew signal output
rlabel metal3 s 198962 29792 199762 29912 6 m_out[19]
port 301 nsew signal output
rlabel metal3 s 198962 2184 199762 2304 6 m_out[1]
port 302 nsew signal output
rlabel metal3 s 198962 31424 199762 31544 6 m_out[20]
port 303 nsew signal output
rlabel metal3 s 198962 32920 199762 33040 6 m_out[21]
port 304 nsew signal output
rlabel metal3 s 198962 34416 199762 34536 6 m_out[22]
port 305 nsew signal output
rlabel metal3 s 198962 36048 199762 36168 6 m_out[23]
port 306 nsew signal output
rlabel metal3 s 198962 37544 199762 37664 6 m_out[24]
port 307 nsew signal output
rlabel metal3 s 198962 39040 199762 39160 6 m_out[25]
port 308 nsew signal output
rlabel metal3 s 198962 40672 199762 40792 6 m_out[26]
port 309 nsew signal output
rlabel metal3 s 198962 42168 199762 42288 6 m_out[27]
port 310 nsew signal output
rlabel metal3 s 198962 43664 199762 43784 6 m_out[28]
port 311 nsew signal output
rlabel metal3 s 198962 45296 199762 45416 6 m_out[29]
port 312 nsew signal output
rlabel metal3 s 198962 3680 199762 3800 6 m_out[2]
port 313 nsew signal output
rlabel metal3 s 198962 46792 199762 46912 6 m_out[30]
port 314 nsew signal output
rlabel metal3 s 198962 48288 199762 48408 6 m_out[31]
port 315 nsew signal output
rlabel metal3 s 198962 49920 199762 50040 6 m_out[32]
port 316 nsew signal output
rlabel metal3 s 198962 51416 199762 51536 6 m_out[33]
port 317 nsew signal output
rlabel metal3 s 198962 52912 199762 53032 6 m_out[34]
port 318 nsew signal output
rlabel metal3 s 198962 54544 199762 54664 6 m_out[35]
port 319 nsew signal output
rlabel metal3 s 198962 56040 199762 56160 6 m_out[36]
port 320 nsew signal output
rlabel metal3 s 198962 57536 199762 57656 6 m_out[37]
port 321 nsew signal output
rlabel metal3 s 198962 59032 199762 59152 6 m_out[38]
port 322 nsew signal output
rlabel metal3 s 198962 60664 199762 60784 6 m_out[39]
port 323 nsew signal output
rlabel metal3 s 198962 5176 199762 5296 6 m_out[3]
port 324 nsew signal output
rlabel metal3 s 198962 62160 199762 62280 6 m_out[40]
port 325 nsew signal output
rlabel metal3 s 198962 63656 199762 63776 6 m_out[41]
port 326 nsew signal output
rlabel metal3 s 198962 65288 199762 65408 6 m_out[42]
port 327 nsew signal output
rlabel metal3 s 198962 66784 199762 66904 6 m_out[43]
port 328 nsew signal output
rlabel metal3 s 198962 68280 199762 68400 6 m_out[44]
port 329 nsew signal output
rlabel metal3 s 198962 69912 199762 70032 6 m_out[45]
port 330 nsew signal output
rlabel metal3 s 198962 71408 199762 71528 6 m_out[46]
port 331 nsew signal output
rlabel metal3 s 198962 72904 199762 73024 6 m_out[47]
port 332 nsew signal output
rlabel metal3 s 198962 74536 199762 74656 6 m_out[48]
port 333 nsew signal output
rlabel metal3 s 198962 76032 199762 76152 6 m_out[49]
port 334 nsew signal output
rlabel metal3 s 198962 6808 199762 6928 6 m_out[4]
port 335 nsew signal output
rlabel metal3 s 198962 77528 199762 77648 6 m_out[50]
port 336 nsew signal output
rlabel metal3 s 198962 79160 199762 79280 6 m_out[51]
port 337 nsew signal output
rlabel metal3 s 198962 80656 199762 80776 6 m_out[52]
port 338 nsew signal output
rlabel metal3 s 198962 82152 199762 82272 6 m_out[53]
port 339 nsew signal output
rlabel metal3 s 198962 83784 199762 83904 6 m_out[54]
port 340 nsew signal output
rlabel metal3 s 198962 85280 199762 85400 6 m_out[55]
port 341 nsew signal output
rlabel metal3 s 198962 86776 199762 86896 6 m_out[56]
port 342 nsew signal output
rlabel metal3 s 198962 88272 199762 88392 6 m_out[57]
port 343 nsew signal output
rlabel metal3 s 198962 89904 199762 90024 6 m_out[58]
port 344 nsew signal output
rlabel metal3 s 198962 91400 199762 91520 6 m_out[59]
port 345 nsew signal output
rlabel metal3 s 198962 8304 199762 8424 6 m_out[5]
port 346 nsew signal output
rlabel metal3 s 198962 92896 199762 93016 6 m_out[60]
port 347 nsew signal output
rlabel metal3 s 198962 94528 199762 94648 6 m_out[61]
port 348 nsew signal output
rlabel metal3 s 198962 96024 199762 96144 6 m_out[62]
port 349 nsew signal output
rlabel metal3 s 198962 97520 199762 97640 6 m_out[63]
port 350 nsew signal output
rlabel metal3 s 198962 99152 199762 99272 6 m_out[64]
port 351 nsew signal output
rlabel metal3 s 198962 100648 199762 100768 6 m_out[65]
port 352 nsew signal output
rlabel metal3 s 198962 102144 199762 102264 6 m_out[66]
port 353 nsew signal output
rlabel metal3 s 198962 103776 199762 103896 6 m_out[67]
port 354 nsew signal output
rlabel metal3 s 198962 105272 199762 105392 6 m_out[68]
port 355 nsew signal output
rlabel metal3 s 198962 106768 199762 106888 6 m_out[69]
port 356 nsew signal output
rlabel metal3 s 198962 9800 199762 9920 6 m_out[6]
port 357 nsew signal output
rlabel metal3 s 198962 108400 199762 108520 6 m_out[70]
port 358 nsew signal output
rlabel metal3 s 198962 109896 199762 110016 6 m_out[71]
port 359 nsew signal output
rlabel metal3 s 198962 111392 199762 111512 6 m_out[72]
port 360 nsew signal output
rlabel metal3 s 198962 113024 199762 113144 6 m_out[73]
port 361 nsew signal output
rlabel metal3 s 198962 114520 199762 114640 6 m_out[74]
port 362 nsew signal output
rlabel metal3 s 198962 116016 199762 116136 6 m_out[75]
port 363 nsew signal output
rlabel metal3 s 198962 117512 199762 117632 6 m_out[76]
port 364 nsew signal output
rlabel metal3 s 198962 119144 199762 119264 6 m_out[77]
port 365 nsew signal output
rlabel metal3 s 198962 120640 199762 120760 6 m_out[78]
port 366 nsew signal output
rlabel metal3 s 198962 122136 199762 122256 6 m_out[79]
port 367 nsew signal output
rlabel metal3 s 198962 11432 199762 11552 6 m_out[7]
port 368 nsew signal output
rlabel metal3 s 198962 123768 199762 123888 6 m_out[80]
port 369 nsew signal output
rlabel metal3 s 198962 125264 199762 125384 6 m_out[81]
port 370 nsew signal output
rlabel metal3 s 198962 126760 199762 126880 6 m_out[82]
port 371 nsew signal output
rlabel metal3 s 198962 128392 199762 128512 6 m_out[83]
port 372 nsew signal output
rlabel metal3 s 198962 129888 199762 130008 6 m_out[84]
port 373 nsew signal output
rlabel metal3 s 198962 131384 199762 131504 6 m_out[85]
port 374 nsew signal output
rlabel metal3 s 198962 133016 199762 133136 6 m_out[86]
port 375 nsew signal output
rlabel metal3 s 198962 134512 199762 134632 6 m_out[87]
port 376 nsew signal output
rlabel metal3 s 198962 136008 199762 136128 6 m_out[88]
port 377 nsew signal output
rlabel metal3 s 198962 137640 199762 137760 6 m_out[89]
port 378 nsew signal output
rlabel metal3 s 198962 12928 199762 13048 6 m_out[8]
port 379 nsew signal output
rlabel metal3 s 198962 139136 199762 139256 6 m_out[90]
port 380 nsew signal output
rlabel metal3 s 198962 140632 199762 140752 6 m_out[91]
port 381 nsew signal output
rlabel metal3 s 198962 142264 199762 142384 6 m_out[92]
port 382 nsew signal output
rlabel metal3 s 198962 143760 199762 143880 6 m_out[93]
port 383 nsew signal output
rlabel metal3 s 198962 145256 199762 145376 6 m_out[94]
port 384 nsew signal output
rlabel metal3 s 198962 146752 199762 146872 6 m_out[95]
port 385 nsew signal output
rlabel metal3 s 198962 148384 199762 148504 6 m_out[96]
port 386 nsew signal output
rlabel metal3 s 198962 149880 199762 150000 6 m_out[97]
port 387 nsew signal output
rlabel metal3 s 198962 151376 199762 151496 6 m_out[98]
port 388 nsew signal output
rlabel metal3 s 198962 153008 199762 153128 6 m_out[99]
port 389 nsew signal output
rlabel metal3 s 198962 14424 199762 14544 6 m_out[9]
port 390 nsew signal output
rlabel metal4 s 188290 2128 188610 197520 6 vccd1
port 391 nsew power bidirectional
rlabel metal4 s 157570 2128 157890 197520 6 vccd1
port 392 nsew power bidirectional
rlabel metal4 s 126850 2128 127170 197520 6 vccd1
port 393 nsew power bidirectional
rlabel metal4 s 96130 2128 96450 197520 6 vccd1
port 394 nsew power bidirectional
rlabel metal4 s 65410 2128 65730 197520 6 vccd1
port 395 nsew power bidirectional
rlabel metal4 s 34690 2128 35010 197520 6 vccd1
port 396 nsew power bidirectional
rlabel metal4 s 3970 2128 4290 197520 6 vccd1
port 397 nsew power bidirectional
rlabel metal4 s 172930 2128 173250 197520 6 vssd1
port 398 nsew ground bidirectional
rlabel metal4 s 142210 2128 142530 197520 6 vssd1
port 399 nsew ground bidirectional
rlabel metal4 s 111490 2128 111810 197520 6 vssd1
port 400 nsew ground bidirectional
rlabel metal4 s 80770 2128 81090 197520 6 vssd1
port 401 nsew ground bidirectional
rlabel metal4 s 50050 2128 50370 197520 6 vssd1
port 402 nsew ground bidirectional
rlabel metal4 s 19330 2128 19650 197520 6 vssd1
port 403 nsew ground bidirectional
rlabel metal4 s 188950 2176 189270 197472 6 vccd2
port 404 nsew power bidirectional
rlabel metal4 s 158230 2176 158550 197472 6 vccd2
port 405 nsew power bidirectional
rlabel metal4 s 127510 2176 127830 197472 6 vccd2
port 406 nsew power bidirectional
rlabel metal4 s 96790 2176 97110 197472 6 vccd2
port 407 nsew power bidirectional
rlabel metal4 s 66070 2176 66390 197472 6 vccd2
port 408 nsew power bidirectional
rlabel metal4 s 35350 2176 35670 197472 6 vccd2
port 409 nsew power bidirectional
rlabel metal4 s 4630 2176 4950 197472 6 vccd2
port 410 nsew power bidirectional
rlabel metal4 s 173590 2176 173910 197472 6 vssd2
port 411 nsew ground bidirectional
rlabel metal4 s 142870 2176 143190 197472 6 vssd2
port 412 nsew ground bidirectional
rlabel metal4 s 112150 2176 112470 197472 6 vssd2
port 413 nsew ground bidirectional
rlabel metal4 s 81430 2176 81750 197472 6 vssd2
port 414 nsew ground bidirectional
rlabel metal4 s 50710 2176 51030 197472 6 vssd2
port 415 nsew ground bidirectional
rlabel metal4 s 19990 2176 20310 197472 6 vssd2
port 416 nsew ground bidirectional
rlabel metal4 s 189610 2176 189930 197472 6 vdda1
port 417 nsew power bidirectional
rlabel metal4 s 158890 2176 159210 197472 6 vdda1
port 418 nsew power bidirectional
rlabel metal4 s 128170 2176 128490 197472 6 vdda1
port 419 nsew power bidirectional
rlabel metal4 s 97450 2176 97770 197472 6 vdda1
port 420 nsew power bidirectional
rlabel metal4 s 66730 2176 67050 197472 6 vdda1
port 421 nsew power bidirectional
rlabel metal4 s 36010 2176 36330 197472 6 vdda1
port 422 nsew power bidirectional
rlabel metal4 s 5290 2176 5610 197472 6 vdda1
port 423 nsew power bidirectional
rlabel metal4 s 174250 2176 174570 197472 6 vssa1
port 424 nsew ground bidirectional
rlabel metal4 s 143530 2176 143850 197472 6 vssa1
port 425 nsew ground bidirectional
rlabel metal4 s 112810 2176 113130 197472 6 vssa1
port 426 nsew ground bidirectional
rlabel metal4 s 82090 2176 82410 197472 6 vssa1
port 427 nsew ground bidirectional
rlabel metal4 s 51370 2176 51690 197472 6 vssa1
port 428 nsew ground bidirectional
rlabel metal4 s 20650 2176 20970 197472 6 vssa1
port 429 nsew ground bidirectional
rlabel metal4 s 190270 2176 190590 197472 6 vdda2
port 430 nsew power bidirectional
rlabel metal4 s 159550 2176 159870 197472 6 vdda2
port 431 nsew power bidirectional
rlabel metal4 s 128830 2176 129150 197472 6 vdda2
port 432 nsew power bidirectional
rlabel metal4 s 98110 2176 98430 197472 6 vdda2
port 433 nsew power bidirectional
rlabel metal4 s 67390 2176 67710 197472 6 vdda2
port 434 nsew power bidirectional
rlabel metal4 s 36670 2176 36990 197472 6 vdda2
port 435 nsew power bidirectional
rlabel metal4 s 5950 2176 6270 197472 6 vdda2
port 436 nsew power bidirectional
rlabel metal4 s 174910 2176 175230 197472 6 vssa2
port 437 nsew ground bidirectional
rlabel metal4 s 144190 2176 144510 197472 6 vssa2
port 438 nsew ground bidirectional
rlabel metal4 s 113470 2176 113790 197472 6 vssa2
port 439 nsew ground bidirectional
rlabel metal4 s 82750 2176 83070 197472 6 vssa2
port 440 nsew ground bidirectional
rlabel metal4 s 52030 2176 52350 197472 6 vssa2
port 441 nsew ground bidirectional
rlabel metal4 s 21310 2176 21630 197472 6 vssa2
port 442 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 199762 200025
string LEFview TRUE
string GDS_FILE /project/openlane/multiply_4/runs/multiply_4/results/magic/multiply_4.gds
string GDS_END 123972538
string GDS_START 399520
<< end >>

