magic
tech sky130A
magscale 1 2
timestamp 1610964531
<< obsli1 >>
rect 1104 655 219391 216113
<< obsm1 >>
rect 14 624 219958 216972
<< metal2 >>
rect 478 217696 534 218496
rect 1490 217696 1546 218496
rect 2502 217696 2558 218496
rect 3514 217696 3570 218496
rect 4526 217696 4582 218496
rect 5538 217696 5594 218496
rect 6550 217696 6606 218496
rect 7562 217696 7618 218496
rect 8574 217696 8630 218496
rect 9586 217696 9642 218496
rect 10598 217696 10654 218496
rect 11610 217696 11666 218496
rect 12622 217696 12678 218496
rect 13634 217696 13690 218496
rect 14646 217696 14702 218496
rect 15658 217696 15714 218496
rect 16670 217696 16726 218496
rect 17682 217696 17738 218496
rect 18694 217696 18750 218496
rect 19706 217696 19762 218496
rect 20718 217696 20774 218496
rect 21730 217696 21786 218496
rect 22742 217696 22798 218496
rect 23754 217696 23810 218496
rect 24766 217696 24822 218496
rect 25778 217696 25834 218496
rect 26790 217696 26846 218496
rect 27802 217696 27858 218496
rect 28814 217696 28870 218496
rect 29826 217696 29882 218496
rect 30838 217696 30894 218496
rect 31850 217696 31906 218496
rect 32862 217696 32918 218496
rect 33874 217696 33930 218496
rect 34886 217696 34942 218496
rect 35898 217696 35954 218496
rect 36910 217696 36966 218496
rect 37922 217696 37978 218496
rect 38934 217696 38990 218496
rect 39946 217696 40002 218496
rect 40958 217696 41014 218496
rect 41970 217696 42026 218496
rect 42982 217696 43038 218496
rect 43994 217696 44050 218496
rect 45006 217696 45062 218496
rect 46018 217696 46074 218496
rect 47030 217696 47086 218496
rect 48042 217696 48098 218496
rect 49054 217696 49110 218496
rect 50066 217696 50122 218496
rect 51078 217696 51134 218496
rect 52090 217696 52146 218496
rect 53102 217696 53158 218496
rect 54114 217696 54170 218496
rect 55126 217696 55182 218496
rect 56230 217696 56286 218496
rect 57242 217696 57298 218496
rect 58254 217696 58310 218496
rect 59266 217696 59322 218496
rect 60278 217696 60334 218496
rect 61290 217696 61346 218496
rect 62302 217696 62358 218496
rect 63314 217696 63370 218496
rect 64326 217696 64382 218496
rect 65338 217696 65394 218496
rect 66350 217696 66406 218496
rect 67362 217696 67418 218496
rect 68374 217696 68430 218496
rect 69386 217696 69442 218496
rect 70398 217696 70454 218496
rect 71410 217696 71466 218496
rect 72422 217696 72478 218496
rect 73434 217696 73490 218496
rect 74446 217696 74502 218496
rect 75458 217696 75514 218496
rect 76470 217696 76526 218496
rect 77482 217696 77538 218496
rect 78494 217696 78550 218496
rect 79506 217696 79562 218496
rect 80518 217696 80574 218496
rect 81530 217696 81586 218496
rect 82542 217696 82598 218496
rect 83554 217696 83610 218496
rect 84566 217696 84622 218496
rect 85578 217696 85634 218496
rect 86590 217696 86646 218496
rect 87602 217696 87658 218496
rect 88614 217696 88670 218496
rect 89626 217696 89682 218496
rect 90638 217696 90694 218496
rect 91650 217696 91706 218496
rect 92662 217696 92718 218496
rect 93674 217696 93730 218496
rect 94686 217696 94742 218496
rect 95698 217696 95754 218496
rect 96710 217696 96766 218496
rect 97722 217696 97778 218496
rect 98734 217696 98790 218496
rect 99746 217696 99802 218496
rect 100758 217696 100814 218496
rect 101770 217696 101826 218496
rect 102782 217696 102838 218496
rect 103794 217696 103850 218496
rect 104806 217696 104862 218496
rect 105818 217696 105874 218496
rect 106830 217696 106886 218496
rect 107842 217696 107898 218496
rect 108854 217696 108910 218496
rect 109866 217696 109922 218496
rect 110970 217696 111026 218496
rect 111982 217696 112038 218496
rect 112994 217696 113050 218496
rect 114006 217696 114062 218496
rect 115018 217696 115074 218496
rect 116030 217696 116086 218496
rect 117042 217696 117098 218496
rect 118054 217696 118110 218496
rect 119066 217696 119122 218496
rect 120078 217696 120134 218496
rect 121090 217696 121146 218496
rect 122102 217696 122158 218496
rect 123114 217696 123170 218496
rect 124126 217696 124182 218496
rect 125138 217696 125194 218496
rect 126150 217696 126206 218496
rect 127162 217696 127218 218496
rect 128174 217696 128230 218496
rect 129186 217696 129242 218496
rect 130198 217696 130254 218496
rect 131210 217696 131266 218496
rect 132222 217696 132278 218496
rect 133234 217696 133290 218496
rect 134246 217696 134302 218496
rect 135258 217696 135314 218496
rect 136270 217696 136326 218496
rect 137282 217696 137338 218496
rect 138294 217696 138350 218496
rect 139306 217696 139362 218496
rect 140318 217696 140374 218496
rect 141330 217696 141386 218496
rect 142342 217696 142398 218496
rect 143354 217696 143410 218496
rect 144366 217696 144422 218496
rect 145378 217696 145434 218496
rect 146390 217696 146446 218496
rect 147402 217696 147458 218496
rect 148414 217696 148470 218496
rect 149426 217696 149482 218496
rect 150438 217696 150494 218496
rect 151450 217696 151506 218496
rect 152462 217696 152518 218496
rect 153474 217696 153530 218496
rect 154486 217696 154542 218496
rect 155498 217696 155554 218496
rect 156510 217696 156566 218496
rect 157522 217696 157578 218496
rect 158534 217696 158590 218496
rect 159546 217696 159602 218496
rect 160558 217696 160614 218496
rect 161570 217696 161626 218496
rect 162582 217696 162638 218496
rect 163594 217696 163650 218496
rect 164606 217696 164662 218496
rect 165710 217696 165766 218496
rect 166722 217696 166778 218496
rect 167734 217696 167790 218496
rect 168746 217696 168802 218496
rect 169758 217696 169814 218496
rect 170770 217696 170826 218496
rect 171782 217696 171838 218496
rect 172794 217696 172850 218496
rect 173806 217696 173862 218496
rect 174818 217696 174874 218496
rect 175830 217696 175886 218496
rect 176842 217696 176898 218496
rect 177854 217696 177910 218496
rect 178866 217696 178922 218496
rect 179878 217696 179934 218496
rect 180890 217696 180946 218496
rect 181902 217696 181958 218496
rect 182914 217696 182970 218496
rect 183926 217696 183982 218496
rect 184938 217696 184994 218496
rect 185950 217696 186006 218496
rect 186962 217696 187018 218496
rect 187974 217696 188030 218496
rect 188986 217696 189042 218496
rect 189998 217696 190054 218496
rect 191010 217696 191066 218496
rect 192022 217696 192078 218496
rect 193034 217696 193090 218496
rect 194046 217696 194102 218496
rect 195058 217696 195114 218496
rect 196070 217696 196126 218496
rect 197082 217696 197138 218496
rect 198094 217696 198150 218496
rect 199106 217696 199162 218496
rect 200118 217696 200174 218496
rect 201130 217696 201186 218496
rect 202142 217696 202198 218496
rect 203154 217696 203210 218496
rect 204166 217696 204222 218496
rect 205178 217696 205234 218496
rect 206190 217696 206246 218496
rect 207202 217696 207258 218496
rect 208214 217696 208270 218496
rect 209226 217696 209282 218496
rect 210238 217696 210294 218496
rect 211250 217696 211306 218496
rect 212262 217696 212318 218496
rect 213274 217696 213330 218496
rect 214286 217696 214342 218496
rect 215298 217696 215354 218496
rect 216310 217696 216366 218496
rect 217322 217696 217378 218496
rect 218334 217696 218390 218496
rect 219346 217696 219402 218496
<< obsm2 >>
rect 18 217640 422 217696
rect 590 217640 1434 217696
rect 1602 217640 2446 217696
rect 2614 217640 3458 217696
rect 3626 217640 4470 217696
rect 4638 217640 5482 217696
rect 5650 217640 6494 217696
rect 6662 217640 7506 217696
rect 7674 217640 8518 217696
rect 8686 217640 9530 217696
rect 9698 217640 10542 217696
rect 10710 217640 11554 217696
rect 11722 217640 12566 217696
rect 12734 217640 13578 217696
rect 13746 217640 14590 217696
rect 14758 217640 15602 217696
rect 15770 217640 16614 217696
rect 16782 217640 17626 217696
rect 17794 217640 18638 217696
rect 18806 217640 19650 217696
rect 19818 217640 20662 217696
rect 20830 217640 21674 217696
rect 21842 217640 22686 217696
rect 22854 217640 23698 217696
rect 23866 217640 24710 217696
rect 24878 217640 25722 217696
rect 25890 217640 26734 217696
rect 26902 217640 27746 217696
rect 27914 217640 28758 217696
rect 28926 217640 29770 217696
rect 29938 217640 30782 217696
rect 30950 217640 31794 217696
rect 31962 217640 32806 217696
rect 32974 217640 33818 217696
rect 33986 217640 34830 217696
rect 34998 217640 35842 217696
rect 36010 217640 36854 217696
rect 37022 217640 37866 217696
rect 38034 217640 38878 217696
rect 39046 217640 39890 217696
rect 40058 217640 40902 217696
rect 41070 217640 41914 217696
rect 42082 217640 42926 217696
rect 43094 217640 43938 217696
rect 44106 217640 44950 217696
rect 45118 217640 45962 217696
rect 46130 217640 46974 217696
rect 47142 217640 47986 217696
rect 48154 217640 48998 217696
rect 49166 217640 50010 217696
rect 50178 217640 51022 217696
rect 51190 217640 52034 217696
rect 52202 217640 53046 217696
rect 53214 217640 54058 217696
rect 54226 217640 55070 217696
rect 55238 217640 56174 217696
rect 56342 217640 57186 217696
rect 57354 217640 58198 217696
rect 58366 217640 59210 217696
rect 59378 217640 60222 217696
rect 60390 217640 61234 217696
rect 61402 217640 62246 217696
rect 62414 217640 63258 217696
rect 63426 217640 64270 217696
rect 64438 217640 65282 217696
rect 65450 217640 66294 217696
rect 66462 217640 67306 217696
rect 67474 217640 68318 217696
rect 68486 217640 69330 217696
rect 69498 217640 70342 217696
rect 70510 217640 71354 217696
rect 71522 217640 72366 217696
rect 72534 217640 73378 217696
rect 73546 217640 74390 217696
rect 74558 217640 75402 217696
rect 75570 217640 76414 217696
rect 76582 217640 77426 217696
rect 77594 217640 78438 217696
rect 78606 217640 79450 217696
rect 79618 217640 80462 217696
rect 80630 217640 81474 217696
rect 81642 217640 82486 217696
rect 82654 217640 83498 217696
rect 83666 217640 84510 217696
rect 84678 217640 85522 217696
rect 85690 217640 86534 217696
rect 86702 217640 87546 217696
rect 87714 217640 88558 217696
rect 88726 217640 89570 217696
rect 89738 217640 90582 217696
rect 90750 217640 91594 217696
rect 91762 217640 92606 217696
rect 92774 217640 93618 217696
rect 93786 217640 94630 217696
rect 94798 217640 95642 217696
rect 95810 217640 96654 217696
rect 96822 217640 97666 217696
rect 97834 217640 98678 217696
rect 98846 217640 99690 217696
rect 99858 217640 100702 217696
rect 100870 217640 101714 217696
rect 101882 217640 102726 217696
rect 102894 217640 103738 217696
rect 103906 217640 104750 217696
rect 104918 217640 105762 217696
rect 105930 217640 106774 217696
rect 106942 217640 107786 217696
rect 107954 217640 108798 217696
rect 108966 217640 109810 217696
rect 109978 217640 110914 217696
rect 111082 217640 111926 217696
rect 112094 217640 112938 217696
rect 113106 217640 113950 217696
rect 114118 217640 114962 217696
rect 115130 217640 115974 217696
rect 116142 217640 116986 217696
rect 117154 217640 117998 217696
rect 118166 217640 119010 217696
rect 119178 217640 120022 217696
rect 120190 217640 121034 217696
rect 121202 217640 122046 217696
rect 122214 217640 123058 217696
rect 123226 217640 124070 217696
rect 124238 217640 125082 217696
rect 125250 217640 126094 217696
rect 126262 217640 127106 217696
rect 127274 217640 128118 217696
rect 128286 217640 129130 217696
rect 129298 217640 130142 217696
rect 130310 217640 131154 217696
rect 131322 217640 132166 217696
rect 132334 217640 133178 217696
rect 133346 217640 134190 217696
rect 134358 217640 135202 217696
rect 135370 217640 136214 217696
rect 136382 217640 137226 217696
rect 137394 217640 138238 217696
rect 138406 217640 139250 217696
rect 139418 217640 140262 217696
rect 140430 217640 141274 217696
rect 141442 217640 142286 217696
rect 142454 217640 143298 217696
rect 143466 217640 144310 217696
rect 144478 217640 145322 217696
rect 145490 217640 146334 217696
rect 146502 217640 147346 217696
rect 147514 217640 148358 217696
rect 148526 217640 149370 217696
rect 149538 217640 150382 217696
rect 150550 217640 151394 217696
rect 151562 217640 152406 217696
rect 152574 217640 153418 217696
rect 153586 217640 154430 217696
rect 154598 217640 155442 217696
rect 155610 217640 156454 217696
rect 156622 217640 157466 217696
rect 157634 217640 158478 217696
rect 158646 217640 159490 217696
rect 159658 217640 160502 217696
rect 160670 217640 161514 217696
rect 161682 217640 162526 217696
rect 162694 217640 163538 217696
rect 163706 217640 164550 217696
rect 164718 217640 165654 217696
rect 165822 217640 166666 217696
rect 166834 217640 167678 217696
rect 167846 217640 168690 217696
rect 168858 217640 169702 217696
rect 169870 217640 170714 217696
rect 170882 217640 171726 217696
rect 171894 217640 172738 217696
rect 172906 217640 173750 217696
rect 173918 217640 174762 217696
rect 174930 217640 175774 217696
rect 175942 217640 176786 217696
rect 176954 217640 177798 217696
rect 177966 217640 178810 217696
rect 178978 217640 179822 217696
rect 179990 217640 180834 217696
rect 181002 217640 181846 217696
rect 182014 217640 182858 217696
rect 183026 217640 183870 217696
rect 184038 217640 184882 217696
rect 185050 217640 185894 217696
rect 186062 217640 186906 217696
rect 187074 217640 187918 217696
rect 188086 217640 188930 217696
rect 189098 217640 189942 217696
rect 190110 217640 190954 217696
rect 191122 217640 191966 217696
rect 192134 217640 192978 217696
rect 193146 217640 193990 217696
rect 194158 217640 195002 217696
rect 195170 217640 196014 217696
rect 196182 217640 197026 217696
rect 197194 217640 198038 217696
rect 198206 217640 199050 217696
rect 199218 217640 200062 217696
rect 200230 217640 201074 217696
rect 201242 217640 202086 217696
rect 202254 217640 203098 217696
rect 203266 217640 204110 217696
rect 204278 217640 205122 217696
rect 205290 217640 206134 217696
rect 206302 217640 207146 217696
rect 207314 217640 208158 217696
rect 208326 217640 209170 217696
rect 209338 217640 210182 217696
rect 210350 217640 211194 217696
rect 211362 217640 212206 217696
rect 212374 217640 213218 217696
rect 213386 217640 214230 217696
rect 214398 217640 215242 217696
rect 215410 217640 216254 217696
rect 216422 217640 217266 217696
rect 217434 217640 218278 217696
rect 218446 217640 219290 217696
rect 219458 217640 219952 217696
rect 18 23 219952 217640
<< metal3 >>
rect 0 216920 800 217040
rect 0 213928 800 214048
rect 0 210800 800 210920
rect 0 207808 800 207928
rect 0 204680 800 204800
rect 0 201688 800 201808
rect 0 198560 800 198680
rect 0 195568 800 195688
rect 0 192440 800 192560
rect 0 189448 800 189568
rect 0 186320 800 186440
rect 0 183328 800 183448
rect 0 180200 800 180320
rect 0 177208 800 177328
rect 0 174080 800 174200
rect 0 171088 800 171208
rect 0 167960 800 168080
rect 0 164968 800 165088
rect 0 161976 800 162096
rect 0 158848 800 158968
rect 0 155856 800 155976
rect 0 152728 800 152848
rect 0 149736 800 149856
rect 0 146608 800 146728
rect 0 143616 800 143736
rect 0 140488 800 140608
rect 0 137496 800 137616
rect 0 134368 800 134488
rect 0 131376 800 131496
rect 0 128248 800 128368
rect 0 125256 800 125376
rect 0 122128 800 122248
rect 0 119136 800 119256
rect 0 116008 800 116128
rect 0 113016 800 113136
rect 0 110024 800 110144
rect 0 106896 800 107016
rect 0 103904 800 104024
rect 0 100776 800 100896
rect 0 97784 800 97904
rect 0 94656 800 94776
rect 0 91664 800 91784
rect 0 88536 800 88656
rect 0 85544 800 85664
rect 0 82416 800 82536
rect 0 79424 800 79544
rect 0 76296 800 76416
rect 0 73304 800 73424
rect 0 70176 800 70296
rect 0 67184 800 67304
rect 0 64056 800 64176
rect 0 61064 800 61184
rect 0 57936 800 58056
rect 0 54944 800 55064
rect 0 51952 800 52072
rect 0 48824 800 48944
rect 0 45832 800 45952
rect 0 42704 800 42824
rect 0 39712 800 39832
rect 0 36584 800 36704
rect 0 33592 800 33712
rect 0 30464 800 30584
rect 0 27472 800 27592
rect 0 24344 800 24464
rect 0 21352 800 21472
rect 0 18224 800 18344
rect 0 15232 800 15352
rect 0 12104 800 12224
rect 0 9112 800 9232
rect 0 5984 800 6104
rect 0 2992 800 3112
rect 0 0 800 120
<< obsm3 >>
rect 13 217120 219867 217149
rect 880 216840 219867 217120
rect 13 214128 219867 216840
rect 880 213848 219867 214128
rect 13 211000 219867 213848
rect 880 210720 219867 211000
rect 13 208008 219867 210720
rect 880 207728 219867 208008
rect 13 204880 219867 207728
rect 880 204600 219867 204880
rect 13 201888 219867 204600
rect 880 201608 219867 201888
rect 13 198760 219867 201608
rect 880 198480 219867 198760
rect 13 195768 219867 198480
rect 880 195488 219867 195768
rect 13 192640 219867 195488
rect 880 192360 219867 192640
rect 13 189648 219867 192360
rect 880 189368 219867 189648
rect 13 186520 219867 189368
rect 880 186240 219867 186520
rect 13 183528 219867 186240
rect 880 183248 219867 183528
rect 13 180400 219867 183248
rect 880 180120 219867 180400
rect 13 177408 219867 180120
rect 880 177128 219867 177408
rect 13 174280 219867 177128
rect 880 174000 219867 174280
rect 13 171288 219867 174000
rect 880 171008 219867 171288
rect 13 168160 219867 171008
rect 880 167880 219867 168160
rect 13 165168 219867 167880
rect 880 164888 219867 165168
rect 13 162176 219867 164888
rect 880 161896 219867 162176
rect 13 159048 219867 161896
rect 880 158768 219867 159048
rect 13 156056 219867 158768
rect 880 155776 219867 156056
rect 13 152928 219867 155776
rect 880 152648 219867 152928
rect 13 149936 219867 152648
rect 880 149656 219867 149936
rect 13 146808 219867 149656
rect 880 146528 219867 146808
rect 13 143816 219867 146528
rect 880 143536 219867 143816
rect 13 140688 219867 143536
rect 880 140408 219867 140688
rect 13 137696 219867 140408
rect 880 137416 219867 137696
rect 13 134568 219867 137416
rect 880 134288 219867 134568
rect 13 131576 219867 134288
rect 880 131296 219867 131576
rect 13 128448 219867 131296
rect 880 128168 219867 128448
rect 13 125456 219867 128168
rect 880 125176 219867 125456
rect 13 122328 219867 125176
rect 880 122048 219867 122328
rect 13 119336 219867 122048
rect 880 119056 219867 119336
rect 13 116208 219867 119056
rect 880 115928 219867 116208
rect 13 113216 219867 115928
rect 880 112936 219867 113216
rect 13 110224 219867 112936
rect 880 109944 219867 110224
rect 13 107096 219867 109944
rect 880 106816 219867 107096
rect 13 104104 219867 106816
rect 880 103824 219867 104104
rect 13 100976 219867 103824
rect 880 100696 219867 100976
rect 13 97984 219867 100696
rect 880 97704 219867 97984
rect 13 94856 219867 97704
rect 880 94576 219867 94856
rect 13 91864 219867 94576
rect 880 91584 219867 91864
rect 13 88736 219867 91584
rect 880 88456 219867 88736
rect 13 85744 219867 88456
rect 880 85464 219867 85744
rect 13 82616 219867 85464
rect 880 82336 219867 82616
rect 13 79624 219867 82336
rect 880 79344 219867 79624
rect 13 76496 219867 79344
rect 880 76216 219867 76496
rect 13 73504 219867 76216
rect 880 73224 219867 73504
rect 13 70376 219867 73224
rect 880 70096 219867 70376
rect 13 67384 219867 70096
rect 880 67104 219867 67384
rect 13 64256 219867 67104
rect 880 63976 219867 64256
rect 13 61264 219867 63976
rect 880 60984 219867 61264
rect 13 58136 219867 60984
rect 880 57856 219867 58136
rect 13 55144 219867 57856
rect 880 54864 219867 55144
rect 13 52152 219867 54864
rect 880 51872 219867 52152
rect 13 49024 219867 51872
rect 880 48744 219867 49024
rect 13 46032 219867 48744
rect 880 45752 219867 46032
rect 13 42904 219867 45752
rect 880 42624 219867 42904
rect 13 39912 219867 42624
rect 880 39632 219867 39912
rect 13 36784 219867 39632
rect 880 36504 219867 36784
rect 13 33792 219867 36504
rect 880 33512 219867 33792
rect 13 30664 219867 33512
rect 880 30384 219867 30664
rect 13 27672 219867 30384
rect 880 27392 219867 27672
rect 13 24544 219867 27392
rect 880 24264 219867 24544
rect 13 21552 219867 24264
rect 880 21272 219867 21552
rect 13 18424 219867 21272
rect 880 18144 219867 18424
rect 13 15432 219867 18144
rect 880 15152 219867 15432
rect 13 12304 219867 15152
rect 880 12024 219867 12304
rect 13 9312 219867 12024
rect 880 9032 219867 9312
rect 13 6184 219867 9032
rect 880 5904 219867 6184
rect 13 3192 219867 5904
rect 880 2912 219867 3192
rect 13 200 219867 2912
rect 880 27 219867 200
<< metal4 >>
rect 4208 624 4528 216144
rect 4868 672 5188 216096
rect 5528 672 5848 216096
rect 6188 672 6508 216096
rect 19568 624 19888 216144
rect 20228 672 20548 216096
rect 20888 672 21208 216096
rect 21548 672 21868 216096
rect 34928 624 35248 216144
rect 35588 672 35908 216096
rect 36248 672 36568 216096
rect 36908 672 37228 216096
rect 50288 624 50608 216144
rect 50948 672 51268 216096
rect 51608 672 51928 216096
rect 52268 672 52588 216096
rect 65648 624 65968 216144
rect 66308 672 66628 216096
rect 66968 672 67288 216096
rect 67628 672 67948 216096
rect 81008 624 81328 216144
rect 81668 672 81988 216096
rect 82328 672 82648 216096
rect 82988 672 83308 216096
rect 96368 624 96688 216144
rect 97028 672 97348 216096
rect 97688 672 98008 216096
rect 98348 672 98668 216096
rect 111728 624 112048 216144
rect 112388 672 112708 216096
rect 113048 672 113368 216096
rect 113708 672 114028 216096
rect 127088 624 127408 216144
rect 127748 672 128068 216096
rect 128408 672 128728 216096
rect 129068 672 129388 216096
rect 142448 624 142768 216144
rect 143108 672 143428 216096
rect 143768 672 144088 216096
rect 144428 672 144748 216096
rect 157808 624 158128 216144
rect 158468 672 158788 216096
rect 159128 672 159448 216096
rect 159788 672 160108 216096
rect 173168 624 173488 216144
rect 173828 672 174148 216096
rect 174488 672 174808 216096
rect 175148 672 175468 216096
rect 188528 624 188848 216144
rect 189188 672 189508 216096
rect 189848 672 190168 216096
rect 190508 672 190828 216096
rect 203888 624 204208 216144
rect 204548 672 204868 216096
rect 205208 672 205528 216096
rect 205868 672 206188 216096
<< obsm4 >>
rect 59 216224 218165 217149
rect 59 9139 4128 216224
rect 4608 216176 19488 216224
rect 4608 9139 4788 216176
rect 5268 9139 5448 216176
rect 5928 9139 6108 216176
rect 6588 9139 19488 216176
rect 19968 216176 34848 216224
rect 19968 9139 20148 216176
rect 20628 9139 20808 216176
rect 21288 9139 21468 216176
rect 21948 9139 34848 216176
rect 35328 216176 50208 216224
rect 35328 9139 35508 216176
rect 35988 9139 36168 216176
rect 36648 9139 36828 216176
rect 37308 9139 50208 216176
rect 50688 216176 65568 216224
rect 50688 9139 50868 216176
rect 51348 9139 51528 216176
rect 52008 9139 52188 216176
rect 52668 9139 65568 216176
rect 66048 216176 80928 216224
rect 66048 9139 66228 216176
rect 66708 9139 66888 216176
rect 67368 9139 67548 216176
rect 68028 9139 80928 216176
rect 81408 216176 96288 216224
rect 81408 9139 81588 216176
rect 82068 9139 82248 216176
rect 82728 9139 82908 216176
rect 83388 9139 96288 216176
rect 96768 216176 111648 216224
rect 96768 9139 96948 216176
rect 97428 9139 97608 216176
rect 98088 9139 98268 216176
rect 98748 9139 111648 216176
rect 112128 216176 127008 216224
rect 112128 9139 112308 216176
rect 112788 9139 112968 216176
rect 113448 9139 113628 216176
rect 114108 9139 127008 216176
rect 127488 216176 142368 216224
rect 127488 9139 127668 216176
rect 128148 9139 128328 216176
rect 128808 9139 128988 216176
rect 129468 9139 142368 216176
rect 142848 216176 157728 216224
rect 142848 9139 143028 216176
rect 143508 9139 143688 216176
rect 144168 9139 144348 216176
rect 144828 9139 157728 216176
rect 158208 216176 173088 216224
rect 158208 9139 158388 216176
rect 158868 9139 159048 216176
rect 159528 9139 159708 216176
rect 160188 9139 173088 216176
rect 173568 216176 188448 216224
rect 173568 9139 173748 216176
rect 174228 9139 174408 216176
rect 174888 9139 175068 216176
rect 175548 9139 188448 216176
rect 188928 216176 203808 216224
rect 188928 9139 189108 216176
rect 189588 9139 189768 216176
rect 190248 9139 190428 216176
rect 190908 9139 203808 216176
rect 204288 216176 218165 216224
rect 204288 9139 204468 216176
rect 204948 9139 205128 216176
rect 205608 9139 205788 216176
rect 206268 9139 218165 216176
<< labels >>
rlabel metal2 s 478 217696 534 218496 6 clk
port 1 nsew signal input
rlabel metal2 s 1490 217696 1546 218496 6 d_in[0]
port 2 nsew signal input
rlabel metal2 s 11610 217696 11666 218496 6 d_in[10]
port 3 nsew signal input
rlabel metal2 s 12622 217696 12678 218496 6 d_in[11]
port 4 nsew signal input
rlabel metal2 s 13634 217696 13690 218496 6 d_in[12]
port 5 nsew signal input
rlabel metal2 s 14646 217696 14702 218496 6 d_in[13]
port 6 nsew signal input
rlabel metal2 s 15658 217696 15714 218496 6 d_in[14]
port 7 nsew signal input
rlabel metal2 s 16670 217696 16726 218496 6 d_in[15]
port 8 nsew signal input
rlabel metal2 s 17682 217696 17738 218496 6 d_in[16]
port 9 nsew signal input
rlabel metal2 s 18694 217696 18750 218496 6 d_in[17]
port 10 nsew signal input
rlabel metal2 s 19706 217696 19762 218496 6 d_in[18]
port 11 nsew signal input
rlabel metal2 s 20718 217696 20774 218496 6 d_in[19]
port 12 nsew signal input
rlabel metal2 s 2502 217696 2558 218496 6 d_in[1]
port 13 nsew signal input
rlabel metal2 s 21730 217696 21786 218496 6 d_in[20]
port 14 nsew signal input
rlabel metal2 s 22742 217696 22798 218496 6 d_in[21]
port 15 nsew signal input
rlabel metal2 s 23754 217696 23810 218496 6 d_in[22]
port 16 nsew signal input
rlabel metal2 s 24766 217696 24822 218496 6 d_in[23]
port 17 nsew signal input
rlabel metal2 s 3514 217696 3570 218496 6 d_in[2]
port 18 nsew signal input
rlabel metal2 s 4526 217696 4582 218496 6 d_in[3]
port 19 nsew signal input
rlabel metal2 s 5538 217696 5594 218496 6 d_in[4]
port 20 nsew signal input
rlabel metal2 s 6550 217696 6606 218496 6 d_in[5]
port 21 nsew signal input
rlabel metal2 s 7562 217696 7618 218496 6 d_in[6]
port 22 nsew signal input
rlabel metal2 s 8574 217696 8630 218496 6 d_in[7]
port 23 nsew signal input
rlabel metal2 s 9586 217696 9642 218496 6 d_in[8]
port 24 nsew signal input
rlabel metal2 s 10598 217696 10654 218496 6 d_in[9]
port 25 nsew signal input
rlabel metal2 s 25778 217696 25834 218496 6 d_out[0]
port 26 nsew signal output
rlabel metal2 s 127162 217696 127218 218496 6 d_out[100]
port 27 nsew signal output
rlabel metal2 s 128174 217696 128230 218496 6 d_out[101]
port 28 nsew signal output
rlabel metal2 s 129186 217696 129242 218496 6 d_out[102]
port 29 nsew signal output
rlabel metal2 s 130198 217696 130254 218496 6 d_out[103]
port 30 nsew signal output
rlabel metal2 s 131210 217696 131266 218496 6 d_out[104]
port 31 nsew signal output
rlabel metal2 s 132222 217696 132278 218496 6 d_out[105]
port 32 nsew signal output
rlabel metal2 s 133234 217696 133290 218496 6 d_out[106]
port 33 nsew signal output
rlabel metal2 s 134246 217696 134302 218496 6 d_out[107]
port 34 nsew signal output
rlabel metal2 s 135258 217696 135314 218496 6 d_out[108]
port 35 nsew signal output
rlabel metal2 s 136270 217696 136326 218496 6 d_out[109]
port 36 nsew signal output
rlabel metal2 s 35898 217696 35954 218496 6 d_out[10]
port 37 nsew signal output
rlabel metal2 s 137282 217696 137338 218496 6 d_out[110]
port 38 nsew signal output
rlabel metal2 s 138294 217696 138350 218496 6 d_out[111]
port 39 nsew signal output
rlabel metal2 s 139306 217696 139362 218496 6 d_out[112]
port 40 nsew signal output
rlabel metal2 s 140318 217696 140374 218496 6 d_out[113]
port 41 nsew signal output
rlabel metal2 s 141330 217696 141386 218496 6 d_out[114]
port 42 nsew signal output
rlabel metal2 s 142342 217696 142398 218496 6 d_out[115]
port 43 nsew signal output
rlabel metal2 s 143354 217696 143410 218496 6 d_out[116]
port 44 nsew signal output
rlabel metal2 s 144366 217696 144422 218496 6 d_out[117]
port 45 nsew signal output
rlabel metal2 s 145378 217696 145434 218496 6 d_out[118]
port 46 nsew signal output
rlabel metal2 s 146390 217696 146446 218496 6 d_out[119]
port 47 nsew signal output
rlabel metal2 s 36910 217696 36966 218496 6 d_out[11]
port 48 nsew signal output
rlabel metal2 s 147402 217696 147458 218496 6 d_out[120]
port 49 nsew signal output
rlabel metal2 s 148414 217696 148470 218496 6 d_out[121]
port 50 nsew signal output
rlabel metal2 s 149426 217696 149482 218496 6 d_out[122]
port 51 nsew signal output
rlabel metal2 s 150438 217696 150494 218496 6 d_out[123]
port 52 nsew signal output
rlabel metal2 s 151450 217696 151506 218496 6 d_out[124]
port 53 nsew signal output
rlabel metal2 s 152462 217696 152518 218496 6 d_out[125]
port 54 nsew signal output
rlabel metal2 s 153474 217696 153530 218496 6 d_out[126]
port 55 nsew signal output
rlabel metal2 s 154486 217696 154542 218496 6 d_out[127]
port 56 nsew signal output
rlabel metal2 s 155498 217696 155554 218496 6 d_out[128]
port 57 nsew signal output
rlabel metal2 s 156510 217696 156566 218496 6 d_out[129]
port 58 nsew signal output
rlabel metal2 s 37922 217696 37978 218496 6 d_out[12]
port 59 nsew signal output
rlabel metal2 s 157522 217696 157578 218496 6 d_out[130]
port 60 nsew signal output
rlabel metal2 s 158534 217696 158590 218496 6 d_out[131]
port 61 nsew signal output
rlabel metal2 s 159546 217696 159602 218496 6 d_out[132]
port 62 nsew signal output
rlabel metal2 s 160558 217696 160614 218496 6 d_out[133]
port 63 nsew signal output
rlabel metal2 s 161570 217696 161626 218496 6 d_out[134]
port 64 nsew signal output
rlabel metal2 s 162582 217696 162638 218496 6 d_out[135]
port 65 nsew signal output
rlabel metal2 s 163594 217696 163650 218496 6 d_out[136]
port 66 nsew signal output
rlabel metal2 s 164606 217696 164662 218496 6 d_out[137]
port 67 nsew signal output
rlabel metal2 s 165710 217696 165766 218496 6 d_out[138]
port 68 nsew signal output
rlabel metal2 s 166722 217696 166778 218496 6 d_out[139]
port 69 nsew signal output
rlabel metal2 s 38934 217696 38990 218496 6 d_out[13]
port 70 nsew signal output
rlabel metal2 s 167734 217696 167790 218496 6 d_out[140]
port 71 nsew signal output
rlabel metal2 s 168746 217696 168802 218496 6 d_out[141]
port 72 nsew signal output
rlabel metal2 s 169758 217696 169814 218496 6 d_out[142]
port 73 nsew signal output
rlabel metal2 s 170770 217696 170826 218496 6 d_out[143]
port 74 nsew signal output
rlabel metal2 s 171782 217696 171838 218496 6 d_out[144]
port 75 nsew signal output
rlabel metal2 s 172794 217696 172850 218496 6 d_out[145]
port 76 nsew signal output
rlabel metal2 s 173806 217696 173862 218496 6 d_out[146]
port 77 nsew signal output
rlabel metal2 s 174818 217696 174874 218496 6 d_out[147]
port 78 nsew signal output
rlabel metal2 s 175830 217696 175886 218496 6 d_out[148]
port 79 nsew signal output
rlabel metal2 s 176842 217696 176898 218496 6 d_out[149]
port 80 nsew signal output
rlabel metal2 s 39946 217696 40002 218496 6 d_out[14]
port 81 nsew signal output
rlabel metal2 s 177854 217696 177910 218496 6 d_out[150]
port 82 nsew signal output
rlabel metal2 s 178866 217696 178922 218496 6 d_out[151]
port 83 nsew signal output
rlabel metal2 s 179878 217696 179934 218496 6 d_out[152]
port 84 nsew signal output
rlabel metal2 s 180890 217696 180946 218496 6 d_out[153]
port 85 nsew signal output
rlabel metal2 s 181902 217696 181958 218496 6 d_out[154]
port 86 nsew signal output
rlabel metal2 s 182914 217696 182970 218496 6 d_out[155]
port 87 nsew signal output
rlabel metal2 s 183926 217696 183982 218496 6 d_out[156]
port 88 nsew signal output
rlabel metal2 s 184938 217696 184994 218496 6 d_out[157]
port 89 nsew signal output
rlabel metal2 s 185950 217696 186006 218496 6 d_out[158]
port 90 nsew signal output
rlabel metal2 s 186962 217696 187018 218496 6 d_out[159]
port 91 nsew signal output
rlabel metal2 s 40958 217696 41014 218496 6 d_out[15]
port 92 nsew signal output
rlabel metal2 s 187974 217696 188030 218496 6 d_out[160]
port 93 nsew signal output
rlabel metal2 s 188986 217696 189042 218496 6 d_out[161]
port 94 nsew signal output
rlabel metal2 s 189998 217696 190054 218496 6 d_out[162]
port 95 nsew signal output
rlabel metal2 s 191010 217696 191066 218496 6 d_out[163]
port 96 nsew signal output
rlabel metal2 s 192022 217696 192078 218496 6 d_out[164]
port 97 nsew signal output
rlabel metal2 s 193034 217696 193090 218496 6 d_out[165]
port 98 nsew signal output
rlabel metal2 s 194046 217696 194102 218496 6 d_out[166]
port 99 nsew signal output
rlabel metal2 s 195058 217696 195114 218496 6 d_out[167]
port 100 nsew signal output
rlabel metal2 s 196070 217696 196126 218496 6 d_out[168]
port 101 nsew signal output
rlabel metal2 s 197082 217696 197138 218496 6 d_out[169]
port 102 nsew signal output
rlabel metal2 s 41970 217696 42026 218496 6 d_out[16]
port 103 nsew signal output
rlabel metal2 s 198094 217696 198150 218496 6 d_out[170]
port 104 nsew signal output
rlabel metal2 s 199106 217696 199162 218496 6 d_out[171]
port 105 nsew signal output
rlabel metal2 s 200118 217696 200174 218496 6 d_out[172]
port 106 nsew signal output
rlabel metal2 s 201130 217696 201186 218496 6 d_out[173]
port 107 nsew signal output
rlabel metal2 s 202142 217696 202198 218496 6 d_out[174]
port 108 nsew signal output
rlabel metal2 s 203154 217696 203210 218496 6 d_out[175]
port 109 nsew signal output
rlabel metal2 s 204166 217696 204222 218496 6 d_out[176]
port 110 nsew signal output
rlabel metal2 s 205178 217696 205234 218496 6 d_out[177]
port 111 nsew signal output
rlabel metal2 s 206190 217696 206246 218496 6 d_out[178]
port 112 nsew signal output
rlabel metal2 s 207202 217696 207258 218496 6 d_out[179]
port 113 nsew signal output
rlabel metal2 s 42982 217696 43038 218496 6 d_out[17]
port 114 nsew signal output
rlabel metal2 s 208214 217696 208270 218496 6 d_out[180]
port 115 nsew signal output
rlabel metal2 s 209226 217696 209282 218496 6 d_out[181]
port 116 nsew signal output
rlabel metal2 s 210238 217696 210294 218496 6 d_out[182]
port 117 nsew signal output
rlabel metal2 s 211250 217696 211306 218496 6 d_out[183]
port 118 nsew signal output
rlabel metal2 s 212262 217696 212318 218496 6 d_out[184]
port 119 nsew signal output
rlabel metal2 s 213274 217696 213330 218496 6 d_out[185]
port 120 nsew signal output
rlabel metal2 s 214286 217696 214342 218496 6 d_out[186]
port 121 nsew signal output
rlabel metal2 s 215298 217696 215354 218496 6 d_out[187]
port 122 nsew signal output
rlabel metal2 s 216310 217696 216366 218496 6 d_out[188]
port 123 nsew signal output
rlabel metal2 s 217322 217696 217378 218496 6 d_out[189]
port 124 nsew signal output
rlabel metal2 s 43994 217696 44050 218496 6 d_out[18]
port 125 nsew signal output
rlabel metal2 s 218334 217696 218390 218496 6 d_out[190]
port 126 nsew signal output
rlabel metal2 s 219346 217696 219402 218496 6 d_out[191]
port 127 nsew signal output
rlabel metal2 s 45006 217696 45062 218496 6 d_out[19]
port 128 nsew signal output
rlabel metal2 s 26790 217696 26846 218496 6 d_out[1]
port 129 nsew signal output
rlabel metal2 s 46018 217696 46074 218496 6 d_out[20]
port 130 nsew signal output
rlabel metal2 s 47030 217696 47086 218496 6 d_out[21]
port 131 nsew signal output
rlabel metal2 s 48042 217696 48098 218496 6 d_out[22]
port 132 nsew signal output
rlabel metal2 s 49054 217696 49110 218496 6 d_out[23]
port 133 nsew signal output
rlabel metal2 s 50066 217696 50122 218496 6 d_out[24]
port 134 nsew signal output
rlabel metal2 s 51078 217696 51134 218496 6 d_out[25]
port 135 nsew signal output
rlabel metal2 s 52090 217696 52146 218496 6 d_out[26]
port 136 nsew signal output
rlabel metal2 s 53102 217696 53158 218496 6 d_out[27]
port 137 nsew signal output
rlabel metal2 s 54114 217696 54170 218496 6 d_out[28]
port 138 nsew signal output
rlabel metal2 s 55126 217696 55182 218496 6 d_out[29]
port 139 nsew signal output
rlabel metal2 s 27802 217696 27858 218496 6 d_out[2]
port 140 nsew signal output
rlabel metal2 s 56230 217696 56286 218496 6 d_out[30]
port 141 nsew signal output
rlabel metal2 s 57242 217696 57298 218496 6 d_out[31]
port 142 nsew signal output
rlabel metal2 s 58254 217696 58310 218496 6 d_out[32]
port 143 nsew signal output
rlabel metal2 s 59266 217696 59322 218496 6 d_out[33]
port 144 nsew signal output
rlabel metal2 s 60278 217696 60334 218496 6 d_out[34]
port 145 nsew signal output
rlabel metal2 s 61290 217696 61346 218496 6 d_out[35]
port 146 nsew signal output
rlabel metal2 s 62302 217696 62358 218496 6 d_out[36]
port 147 nsew signal output
rlabel metal2 s 63314 217696 63370 218496 6 d_out[37]
port 148 nsew signal output
rlabel metal2 s 64326 217696 64382 218496 6 d_out[38]
port 149 nsew signal output
rlabel metal2 s 65338 217696 65394 218496 6 d_out[39]
port 150 nsew signal output
rlabel metal2 s 28814 217696 28870 218496 6 d_out[3]
port 151 nsew signal output
rlabel metal2 s 66350 217696 66406 218496 6 d_out[40]
port 152 nsew signal output
rlabel metal2 s 67362 217696 67418 218496 6 d_out[41]
port 153 nsew signal output
rlabel metal2 s 68374 217696 68430 218496 6 d_out[42]
port 154 nsew signal output
rlabel metal2 s 69386 217696 69442 218496 6 d_out[43]
port 155 nsew signal output
rlabel metal2 s 70398 217696 70454 218496 6 d_out[44]
port 156 nsew signal output
rlabel metal2 s 71410 217696 71466 218496 6 d_out[45]
port 157 nsew signal output
rlabel metal2 s 72422 217696 72478 218496 6 d_out[46]
port 158 nsew signal output
rlabel metal2 s 73434 217696 73490 218496 6 d_out[47]
port 159 nsew signal output
rlabel metal2 s 74446 217696 74502 218496 6 d_out[48]
port 160 nsew signal output
rlabel metal2 s 75458 217696 75514 218496 6 d_out[49]
port 161 nsew signal output
rlabel metal2 s 29826 217696 29882 218496 6 d_out[4]
port 162 nsew signal output
rlabel metal2 s 76470 217696 76526 218496 6 d_out[50]
port 163 nsew signal output
rlabel metal2 s 77482 217696 77538 218496 6 d_out[51]
port 164 nsew signal output
rlabel metal2 s 78494 217696 78550 218496 6 d_out[52]
port 165 nsew signal output
rlabel metal2 s 79506 217696 79562 218496 6 d_out[53]
port 166 nsew signal output
rlabel metal2 s 80518 217696 80574 218496 6 d_out[54]
port 167 nsew signal output
rlabel metal2 s 81530 217696 81586 218496 6 d_out[55]
port 168 nsew signal output
rlabel metal2 s 82542 217696 82598 218496 6 d_out[56]
port 169 nsew signal output
rlabel metal2 s 83554 217696 83610 218496 6 d_out[57]
port 170 nsew signal output
rlabel metal2 s 84566 217696 84622 218496 6 d_out[58]
port 171 nsew signal output
rlabel metal2 s 85578 217696 85634 218496 6 d_out[59]
port 172 nsew signal output
rlabel metal2 s 30838 217696 30894 218496 6 d_out[5]
port 173 nsew signal output
rlabel metal2 s 86590 217696 86646 218496 6 d_out[60]
port 174 nsew signal output
rlabel metal2 s 87602 217696 87658 218496 6 d_out[61]
port 175 nsew signal output
rlabel metal2 s 88614 217696 88670 218496 6 d_out[62]
port 176 nsew signal output
rlabel metal2 s 89626 217696 89682 218496 6 d_out[63]
port 177 nsew signal output
rlabel metal2 s 90638 217696 90694 218496 6 d_out[64]
port 178 nsew signal output
rlabel metal2 s 91650 217696 91706 218496 6 d_out[65]
port 179 nsew signal output
rlabel metal2 s 92662 217696 92718 218496 6 d_out[66]
port 180 nsew signal output
rlabel metal2 s 93674 217696 93730 218496 6 d_out[67]
port 181 nsew signal output
rlabel metal2 s 94686 217696 94742 218496 6 d_out[68]
port 182 nsew signal output
rlabel metal2 s 95698 217696 95754 218496 6 d_out[69]
port 183 nsew signal output
rlabel metal2 s 31850 217696 31906 218496 6 d_out[6]
port 184 nsew signal output
rlabel metal2 s 96710 217696 96766 218496 6 d_out[70]
port 185 nsew signal output
rlabel metal2 s 97722 217696 97778 218496 6 d_out[71]
port 186 nsew signal output
rlabel metal2 s 98734 217696 98790 218496 6 d_out[72]
port 187 nsew signal output
rlabel metal2 s 99746 217696 99802 218496 6 d_out[73]
port 188 nsew signal output
rlabel metal2 s 100758 217696 100814 218496 6 d_out[74]
port 189 nsew signal output
rlabel metal2 s 101770 217696 101826 218496 6 d_out[75]
port 190 nsew signal output
rlabel metal2 s 102782 217696 102838 218496 6 d_out[76]
port 191 nsew signal output
rlabel metal2 s 103794 217696 103850 218496 6 d_out[77]
port 192 nsew signal output
rlabel metal2 s 104806 217696 104862 218496 6 d_out[78]
port 193 nsew signal output
rlabel metal2 s 105818 217696 105874 218496 6 d_out[79]
port 194 nsew signal output
rlabel metal2 s 32862 217696 32918 218496 6 d_out[7]
port 195 nsew signal output
rlabel metal2 s 106830 217696 106886 218496 6 d_out[80]
port 196 nsew signal output
rlabel metal2 s 107842 217696 107898 218496 6 d_out[81]
port 197 nsew signal output
rlabel metal2 s 108854 217696 108910 218496 6 d_out[82]
port 198 nsew signal output
rlabel metal2 s 109866 217696 109922 218496 6 d_out[83]
port 199 nsew signal output
rlabel metal2 s 110970 217696 111026 218496 6 d_out[84]
port 200 nsew signal output
rlabel metal2 s 111982 217696 112038 218496 6 d_out[85]
port 201 nsew signal output
rlabel metal2 s 112994 217696 113050 218496 6 d_out[86]
port 202 nsew signal output
rlabel metal2 s 114006 217696 114062 218496 6 d_out[87]
port 203 nsew signal output
rlabel metal2 s 115018 217696 115074 218496 6 d_out[88]
port 204 nsew signal output
rlabel metal2 s 116030 217696 116086 218496 6 d_out[89]
port 205 nsew signal output
rlabel metal2 s 33874 217696 33930 218496 6 d_out[8]
port 206 nsew signal output
rlabel metal2 s 117042 217696 117098 218496 6 d_out[90]
port 207 nsew signal output
rlabel metal2 s 118054 217696 118110 218496 6 d_out[91]
port 208 nsew signal output
rlabel metal2 s 119066 217696 119122 218496 6 d_out[92]
port 209 nsew signal output
rlabel metal2 s 120078 217696 120134 218496 6 d_out[93]
port 210 nsew signal output
rlabel metal2 s 121090 217696 121146 218496 6 d_out[94]
port 211 nsew signal output
rlabel metal2 s 122102 217696 122158 218496 6 d_out[95]
port 212 nsew signal output
rlabel metal2 s 123114 217696 123170 218496 6 d_out[96]
port 213 nsew signal output
rlabel metal2 s 124126 217696 124182 218496 6 d_out[97]
port 214 nsew signal output
rlabel metal2 s 125138 217696 125194 218496 6 d_out[98]
port 215 nsew signal output
rlabel metal2 s 126150 217696 126206 218496 6 d_out[99]
port 216 nsew signal output
rlabel metal2 s 34886 217696 34942 218496 6 d_out[9]
port 217 nsew signal output
rlabel metal3 s 0 0 800 120 6 w_in[0]
port 218 nsew signal input
rlabel metal3 s 0 30464 800 30584 6 w_in[10]
port 219 nsew signal input
rlabel metal3 s 0 33592 800 33712 6 w_in[11]
port 220 nsew signal input
rlabel metal3 s 0 36584 800 36704 6 w_in[12]
port 221 nsew signal input
rlabel metal3 s 0 39712 800 39832 6 w_in[13]
port 222 nsew signal input
rlabel metal3 s 0 42704 800 42824 6 w_in[14]
port 223 nsew signal input
rlabel metal3 s 0 45832 800 45952 6 w_in[15]
port 224 nsew signal input
rlabel metal3 s 0 48824 800 48944 6 w_in[16]
port 225 nsew signal input
rlabel metal3 s 0 51952 800 52072 6 w_in[17]
port 226 nsew signal input
rlabel metal3 s 0 54944 800 55064 6 w_in[18]
port 227 nsew signal input
rlabel metal3 s 0 57936 800 58056 6 w_in[19]
port 228 nsew signal input
rlabel metal3 s 0 2992 800 3112 6 w_in[1]
port 229 nsew signal input
rlabel metal3 s 0 61064 800 61184 6 w_in[20]
port 230 nsew signal input
rlabel metal3 s 0 64056 800 64176 6 w_in[21]
port 231 nsew signal input
rlabel metal3 s 0 67184 800 67304 6 w_in[22]
port 232 nsew signal input
rlabel metal3 s 0 70176 800 70296 6 w_in[23]
port 233 nsew signal input
rlabel metal3 s 0 73304 800 73424 6 w_in[24]
port 234 nsew signal input
rlabel metal3 s 0 76296 800 76416 6 w_in[25]
port 235 nsew signal input
rlabel metal3 s 0 79424 800 79544 6 w_in[26]
port 236 nsew signal input
rlabel metal3 s 0 82416 800 82536 6 w_in[27]
port 237 nsew signal input
rlabel metal3 s 0 85544 800 85664 6 w_in[28]
port 238 nsew signal input
rlabel metal3 s 0 88536 800 88656 6 w_in[29]
port 239 nsew signal input
rlabel metal3 s 0 5984 800 6104 6 w_in[2]
port 240 nsew signal input
rlabel metal3 s 0 91664 800 91784 6 w_in[30]
port 241 nsew signal input
rlabel metal3 s 0 94656 800 94776 6 w_in[31]
port 242 nsew signal input
rlabel metal3 s 0 97784 800 97904 6 w_in[32]
port 243 nsew signal input
rlabel metal3 s 0 100776 800 100896 6 w_in[33]
port 244 nsew signal input
rlabel metal3 s 0 103904 800 104024 6 w_in[34]
port 245 nsew signal input
rlabel metal3 s 0 106896 800 107016 6 w_in[35]
port 246 nsew signal input
rlabel metal3 s 0 110024 800 110144 6 w_in[36]
port 247 nsew signal input
rlabel metal3 s 0 113016 800 113136 6 w_in[37]
port 248 nsew signal input
rlabel metal3 s 0 116008 800 116128 6 w_in[38]
port 249 nsew signal input
rlabel metal3 s 0 119136 800 119256 6 w_in[39]
port 250 nsew signal input
rlabel metal3 s 0 9112 800 9232 6 w_in[3]
port 251 nsew signal input
rlabel metal3 s 0 122128 800 122248 6 w_in[40]
port 252 nsew signal input
rlabel metal3 s 0 125256 800 125376 6 w_in[41]
port 253 nsew signal input
rlabel metal3 s 0 128248 800 128368 6 w_in[42]
port 254 nsew signal input
rlabel metal3 s 0 131376 800 131496 6 w_in[43]
port 255 nsew signal input
rlabel metal3 s 0 134368 800 134488 6 w_in[44]
port 256 nsew signal input
rlabel metal3 s 0 137496 800 137616 6 w_in[45]
port 257 nsew signal input
rlabel metal3 s 0 140488 800 140608 6 w_in[46]
port 258 nsew signal input
rlabel metal3 s 0 143616 800 143736 6 w_in[47]
port 259 nsew signal input
rlabel metal3 s 0 146608 800 146728 6 w_in[48]
port 260 nsew signal input
rlabel metal3 s 0 149736 800 149856 6 w_in[49]
port 261 nsew signal input
rlabel metal3 s 0 12104 800 12224 6 w_in[4]
port 262 nsew signal input
rlabel metal3 s 0 152728 800 152848 6 w_in[50]
port 263 nsew signal input
rlabel metal3 s 0 155856 800 155976 6 w_in[51]
port 264 nsew signal input
rlabel metal3 s 0 158848 800 158968 6 w_in[52]
port 265 nsew signal input
rlabel metal3 s 0 161976 800 162096 6 w_in[53]
port 266 nsew signal input
rlabel metal3 s 0 164968 800 165088 6 w_in[54]
port 267 nsew signal input
rlabel metal3 s 0 167960 800 168080 6 w_in[55]
port 268 nsew signal input
rlabel metal3 s 0 171088 800 171208 6 w_in[56]
port 269 nsew signal input
rlabel metal3 s 0 174080 800 174200 6 w_in[57]
port 270 nsew signal input
rlabel metal3 s 0 177208 800 177328 6 w_in[58]
port 271 nsew signal input
rlabel metal3 s 0 180200 800 180320 6 w_in[59]
port 272 nsew signal input
rlabel metal3 s 0 15232 800 15352 6 w_in[5]
port 273 nsew signal input
rlabel metal3 s 0 183328 800 183448 6 w_in[60]
port 274 nsew signal input
rlabel metal3 s 0 186320 800 186440 6 w_in[61]
port 275 nsew signal input
rlabel metal3 s 0 189448 800 189568 6 w_in[62]
port 276 nsew signal input
rlabel metal3 s 0 192440 800 192560 6 w_in[63]
port 277 nsew signal input
rlabel metal3 s 0 195568 800 195688 6 w_in[64]
port 278 nsew signal input
rlabel metal3 s 0 198560 800 198680 6 w_in[65]
port 279 nsew signal input
rlabel metal3 s 0 201688 800 201808 6 w_in[66]
port 280 nsew signal input
rlabel metal3 s 0 204680 800 204800 6 w_in[67]
port 281 nsew signal input
rlabel metal3 s 0 207808 800 207928 6 w_in[68]
port 282 nsew signal input
rlabel metal3 s 0 210800 800 210920 6 w_in[69]
port 283 nsew signal input
rlabel metal3 s 0 18224 800 18344 6 w_in[6]
port 284 nsew signal input
rlabel metal3 s 0 213928 800 214048 6 w_in[70]
port 285 nsew signal input
rlabel metal3 s 0 216920 800 217040 6 w_in[71]
port 286 nsew signal input
rlabel metal3 s 0 21352 800 21472 6 w_in[7]
port 287 nsew signal input
rlabel metal3 s 0 24344 800 24464 6 w_in[8]
port 288 nsew signal input
rlabel metal3 s 0 27472 800 27592 6 w_in[9]
port 289 nsew signal input
rlabel metal4 s 188528 624 188848 216144 6 vccd1
port 290 nsew power bidirectional
rlabel metal4 s 157808 624 158128 216144 6 vccd1
port 291 nsew power bidirectional
rlabel metal4 s 127088 624 127408 216144 6 vccd1
port 292 nsew power bidirectional
rlabel metal4 s 96368 624 96688 216144 6 vccd1
port 293 nsew power bidirectional
rlabel metal4 s 65648 624 65968 216144 6 vccd1
port 294 nsew power bidirectional
rlabel metal4 s 34928 624 35248 216144 6 vccd1
port 295 nsew power bidirectional
rlabel metal4 s 4208 624 4528 216144 6 vccd1
port 296 nsew power bidirectional
rlabel metal4 s 203888 624 204208 216144 6 vssd1
port 297 nsew ground bidirectional
rlabel metal4 s 173168 624 173488 216144 6 vssd1
port 298 nsew ground bidirectional
rlabel metal4 s 142448 624 142768 216144 6 vssd1
port 299 nsew ground bidirectional
rlabel metal4 s 111728 624 112048 216144 6 vssd1
port 300 nsew ground bidirectional
rlabel metal4 s 81008 624 81328 216144 6 vssd1
port 301 nsew ground bidirectional
rlabel metal4 s 50288 624 50608 216144 6 vssd1
port 302 nsew ground bidirectional
rlabel metal4 s 19568 624 19888 216144 6 vssd1
port 303 nsew ground bidirectional
rlabel metal4 s 189188 672 189508 216096 6 vccd2
port 304 nsew power bidirectional
rlabel metal4 s 158468 672 158788 216096 6 vccd2
port 305 nsew power bidirectional
rlabel metal4 s 127748 672 128068 216096 6 vccd2
port 306 nsew power bidirectional
rlabel metal4 s 97028 672 97348 216096 6 vccd2
port 307 nsew power bidirectional
rlabel metal4 s 66308 672 66628 216096 6 vccd2
port 308 nsew power bidirectional
rlabel metal4 s 35588 672 35908 216096 6 vccd2
port 309 nsew power bidirectional
rlabel metal4 s 4868 672 5188 216096 6 vccd2
port 310 nsew power bidirectional
rlabel metal4 s 204548 672 204868 216096 6 vssd2
port 311 nsew ground bidirectional
rlabel metal4 s 173828 672 174148 216096 6 vssd2
port 312 nsew ground bidirectional
rlabel metal4 s 143108 672 143428 216096 6 vssd2
port 313 nsew ground bidirectional
rlabel metal4 s 112388 672 112708 216096 6 vssd2
port 314 nsew ground bidirectional
rlabel metal4 s 81668 672 81988 216096 6 vssd2
port 315 nsew ground bidirectional
rlabel metal4 s 50948 672 51268 216096 6 vssd2
port 316 nsew ground bidirectional
rlabel metal4 s 20228 672 20548 216096 6 vssd2
port 317 nsew ground bidirectional
rlabel metal4 s 189848 672 190168 216096 6 vdda1
port 318 nsew power bidirectional
rlabel metal4 s 159128 672 159448 216096 6 vdda1
port 319 nsew power bidirectional
rlabel metal4 s 128408 672 128728 216096 6 vdda1
port 320 nsew power bidirectional
rlabel metal4 s 97688 672 98008 216096 6 vdda1
port 321 nsew power bidirectional
rlabel metal4 s 66968 672 67288 216096 6 vdda1
port 322 nsew power bidirectional
rlabel metal4 s 36248 672 36568 216096 6 vdda1
port 323 nsew power bidirectional
rlabel metal4 s 5528 672 5848 216096 6 vdda1
port 324 nsew power bidirectional
rlabel metal4 s 205208 672 205528 216096 6 vssa1
port 325 nsew ground bidirectional
rlabel metal4 s 174488 672 174808 216096 6 vssa1
port 326 nsew ground bidirectional
rlabel metal4 s 143768 672 144088 216096 6 vssa1
port 327 nsew ground bidirectional
rlabel metal4 s 113048 672 113368 216096 6 vssa1
port 328 nsew ground bidirectional
rlabel metal4 s 82328 672 82648 216096 6 vssa1
port 329 nsew ground bidirectional
rlabel metal4 s 51608 672 51928 216096 6 vssa1
port 330 nsew ground bidirectional
rlabel metal4 s 20888 672 21208 216096 6 vssa1
port 331 nsew ground bidirectional
rlabel metal4 s 190508 672 190828 216096 6 vdda2
port 332 nsew power bidirectional
rlabel metal4 s 159788 672 160108 216096 6 vdda2
port 333 nsew power bidirectional
rlabel metal4 s 129068 672 129388 216096 6 vdda2
port 334 nsew power bidirectional
rlabel metal4 s 98348 672 98668 216096 6 vdda2
port 335 nsew power bidirectional
rlabel metal4 s 67628 672 67948 216096 6 vdda2
port 336 nsew power bidirectional
rlabel metal4 s 36908 672 37228 216096 6 vdda2
port 337 nsew power bidirectional
rlabel metal4 s 6188 672 6508 216096 6 vdda2
port 338 nsew power bidirectional
rlabel metal4 s 205868 672 206188 216096 6 vssa2
port 339 nsew ground bidirectional
rlabel metal4 s 175148 672 175468 216096 6 vssa2
port 340 nsew ground bidirectional
rlabel metal4 s 144428 672 144748 216096 6 vssa2
port 341 nsew ground bidirectional
rlabel metal4 s 113708 672 114028 216096 6 vssa2
port 342 nsew ground bidirectional
rlabel metal4 s 82988 672 83308 216096 6 vssa2
port 343 nsew ground bidirectional
rlabel metal4 s 52268 672 52588 216096 6 vssa2
port 344 nsew ground bidirectional
rlabel metal4 s 21548 672 21868 216096 6 vssa2
port 345 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 219958 218496
string LEFview TRUE
string GDS_FILE /project/openlane/register_file/runs/register_file/results/magic/register_file.gds
string GDS_END 137815432
string GDS_START 221676
<< end >>

