VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dcache
  CLASS BLOCK ;
  FOREIGN dcache ;
  ORIGIN 0.000 0.000 ;
  SIZE 747.890 BY 750.030 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END clk
  PIN d_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END d_in[0]
  PIN d_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END d_in[100]
  PIN d_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END d_in[101]
  PIN d_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 4.000 ;
    END
  END d_in[102]
  PIN d_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END d_in[103]
  PIN d_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 0.000 372.970 4.000 ;
    END
  END d_in[104]
  PIN d_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END d_in[105]
  PIN d_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 0.000 379.870 4.000 ;
    END
  END d_in[106]
  PIN d_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END d_in[107]
  PIN d_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END d_in[108]
  PIN d_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 0.000 390.450 4.000 ;
    END
  END d_in[109]
  PIN d_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END d_in[10]
  PIN d_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END d_in[110]
  PIN d_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 0.000 397.810 4.000 ;
    END
  END d_in[111]
  PIN d_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.750 0.000 401.030 4.000 ;
    END
  END d_in[112]
  PIN d_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END d_in[113]
  PIN d_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END d_in[114]
  PIN d_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 4.000 ;
    END
  END d_in[115]
  PIN d_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.010 0.000 415.290 4.000 ;
    END
  END d_in[116]
  PIN d_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END d_in[117]
  PIN d_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END d_in[118]
  PIN d_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 0.000 425.870 4.000 ;
    END
  END d_in[119]
  PIN d_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END d_in[11]
  PIN d_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 0.000 429.550 4.000 ;
    END
  END d_in[120]
  PIN d_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 4.000 ;
    END
  END d_in[121]
  PIN d_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 4.000 ;
    END
  END d_in[122]
  PIN d_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 0.000 440.130 4.000 ;
    END
  END d_in[123]
  PIN d_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 0.000 443.810 4.000 ;
    END
  END d_in[124]
  PIN d_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END d_in[125]
  PIN d_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 0.000 450.710 4.000 ;
    END
  END d_in[126]
  PIN d_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END d_in[127]
  PIN d_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END d_in[128]
  PIN d_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END d_in[129]
  PIN d_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END d_in[12]
  PIN d_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 0.000 464.970 4.000 ;
    END
  END d_in[130]
  PIN d_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 0.000 468.190 4.000 ;
    END
  END d_in[131]
  PIN d_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END d_in[132]
  PIN d_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 0.000 475.550 4.000 ;
    END
  END d_in[133]
  PIN d_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 0.000 478.770 4.000 ;
    END
  END d_in[134]
  PIN d_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END d_in[135]
  PIN d_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END d_in[136]
  PIN d_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END d_in[137]
  PIN d_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END d_in[138]
  PIN d_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END d_in[139]
  PIN d_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END d_in[13]
  PIN d_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.110 0.000 500.390 4.000 ;
    END
  END d_in[140]
  PIN d_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 0.000 503.610 4.000 ;
    END
  END d_in[141]
  PIN d_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.010 0.000 507.290 4.000 ;
    END
  END d_in[142]
  PIN d_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END d_in[14]
  PIN d_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END d_in[15]
  PIN d_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END d_in[16]
  PIN d_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END d_in[17]
  PIN d_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END d_in[18]
  PIN d_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END d_in[19]
  PIN d_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END d_in[1]
  PIN d_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END d_in[20]
  PIN d_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END d_in[21]
  PIN d_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END d_in[22]
  PIN d_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END d_in[23]
  PIN d_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END d_in[24]
  PIN d_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END d_in[25]
  PIN d_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END d_in[26]
  PIN d_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END d_in[27]
  PIN d_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END d_in[28]
  PIN d_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END d_in[29]
  PIN d_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END d_in[2]
  PIN d_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END d_in[30]
  PIN d_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END d_in[31]
  PIN d_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END d_in[32]
  PIN d_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END d_in[33]
  PIN d_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END d_in[34]
  PIN d_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 4.000 ;
    END
  END d_in[35]
  PIN d_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END d_in[36]
  PIN d_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END d_in[37]
  PIN d_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END d_in[38]
  PIN d_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END d_in[39]
  PIN d_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END d_in[3]
  PIN d_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END d_in[40]
  PIN d_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END d_in[41]
  PIN d_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 4.000 ;
    END
  END d_in[42]
  PIN d_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END d_in[43]
  PIN d_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END d_in[44]
  PIN d_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END d_in[45]
  PIN d_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END d_in[46]
  PIN d_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END d_in[47]
  PIN d_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END d_in[48]
  PIN d_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END d_in[49]
  PIN d_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END d_in[4]
  PIN d_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END d_in[50]
  PIN d_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END d_in[51]
  PIN d_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END d_in[52]
  PIN d_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END d_in[53]
  PIN d_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END d_in[54]
  PIN d_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END d_in[55]
  PIN d_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END d_in[56]
  PIN d_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END d_in[57]
  PIN d_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END d_in[58]
  PIN d_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END d_in[59]
  PIN d_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END d_in[5]
  PIN d_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END d_in[60]
  PIN d_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 0.000 220.710 4.000 ;
    END
  END d_in[61]
  PIN d_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END d_in[62]
  PIN d_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END d_in[63]
  PIN d_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END d_in[64]
  PIN d_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END d_in[65]
  PIN d_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END d_in[66]
  PIN d_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END d_in[67]
  PIN d_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END d_in[68]
  PIN d_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END d_in[69]
  PIN d_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END d_in[6]
  PIN d_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END d_in[70]
  PIN d_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END d_in[71]
  PIN d_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END d_in[72]
  PIN d_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END d_in[73]
  PIN d_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END d_in[74]
  PIN d_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END d_in[75]
  PIN d_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END d_in[76]
  PIN d_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END d_in[77]
  PIN d_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END d_in[78]
  PIN d_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END d_in[79]
  PIN d_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END d_in[7]
  PIN d_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END d_in[80]
  PIN d_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 4.000 ;
    END
  END d_in[81]
  PIN d_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END d_in[82]
  PIN d_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END d_in[83]
  PIN d_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END d_in[84]
  PIN d_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 4.000 ;
    END
  END d_in[85]
  PIN d_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END d_in[86]
  PIN d_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END d_in[87]
  PIN d_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END d_in[88]
  PIN d_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END d_in[89]
  PIN d_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END d_in[8]
  PIN d_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END d_in[90]
  PIN d_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END d_in[91]
  PIN d_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END d_in[92]
  PIN d_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END d_in[93]
  PIN d_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END d_in[94]
  PIN d_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 4.000 ;
    END
  END d_in[95]
  PIN d_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END d_in[96]
  PIN d_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END d_in[97]
  PIN d_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END d_in[98]
  PIN d_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END d_in[99]
  PIN d_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END d_in[9]
  PIN d_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 0.000 510.970 4.000 ;
    END
  END d_out[0]
  PIN d_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 0.000 546.390 4.000 ;
    END
  END d_out[10]
  PIN d_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 0.000 549.610 4.000 ;
    END
  END d_out[11]
  PIN d_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 0.000 553.290 4.000 ;
    END
  END d_out[12]
  PIN d_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END d_out[13]
  PIN d_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 0.000 560.190 4.000 ;
    END
  END d_out[14]
  PIN d_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END d_out[15]
  PIN d_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 0.000 567.550 4.000 ;
    END
  END d_out[16]
  PIN d_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 0.000 570.770 4.000 ;
    END
  END d_out[17]
  PIN d_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 0.000 574.450 4.000 ;
    END
  END d_out[18]
  PIN d_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 0.000 578.130 4.000 ;
    END
  END d_out[19]
  PIN d_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 0.000 514.190 4.000 ;
    END
  END d_out[1]
  PIN d_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 0.000 581.350 4.000 ;
    END
  END d_out[20]
  PIN d_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.750 0.000 585.030 4.000 ;
    END
  END d_out[21]
  PIN d_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.430 0.000 588.710 4.000 ;
    END
  END d_out[22]
  PIN d_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 0.000 592.390 4.000 ;
    END
  END d_out[23]
  PIN d_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 4.000 ;
    END
  END d_out[24]
  PIN d_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END d_out[25]
  PIN d_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.690 0.000 602.970 4.000 ;
    END
  END d_out[26]
  PIN d_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 0.000 606.190 4.000 ;
    END
  END d_out[27]
  PIN d_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 0.000 609.870 4.000 ;
    END
  END d_out[28]
  PIN d_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 0.000 613.550 4.000 ;
    END
  END d_out[29]
  PIN d_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 0.000 517.870 4.000 ;
    END
  END d_out[2]
  PIN d_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.490 0.000 616.770 4.000 ;
    END
  END d_out[30]
  PIN d_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.170 0.000 620.450 4.000 ;
    END
  END d_out[31]
  PIN d_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 0.000 624.130 4.000 ;
    END
  END d_out[32]
  PIN d_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.070 0.000 627.350 4.000 ;
    END
  END d_out[33]
  PIN d_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.750 0.000 631.030 4.000 ;
    END
  END d_out[34]
  PIN d_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 0.000 634.710 4.000 ;
    END
  END d_out[35]
  PIN d_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END d_out[36]
  PIN d_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 0.000 641.610 4.000 ;
    END
  END d_out[37]
  PIN d_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.010 0.000 645.290 4.000 ;
    END
  END d_out[38]
  PIN d_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 0.000 648.970 4.000 ;
    END
  END d_out[39]
  PIN d_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 0.000 521.550 4.000 ;
    END
  END d_out[3]
  PIN d_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.910 0.000 652.190 4.000 ;
    END
  END d_out[40]
  PIN d_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.590 0.000 655.870 4.000 ;
    END
  END d_out[41]
  PIN d_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.270 0.000 659.550 4.000 ;
    END
  END d_out[42]
  PIN d_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 0.000 662.770 4.000 ;
    END
  END d_out[43]
  PIN d_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.170 0.000 666.450 4.000 ;
    END
  END d_out[44]
  PIN d_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END d_out[45]
  PIN d_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END d_out[46]
  PIN d_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 0.000 677.030 4.000 ;
    END
  END d_out[47]
  PIN d_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 0.000 680.710 4.000 ;
    END
  END d_out[48]
  PIN d_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.650 0.000 683.930 4.000 ;
    END
  END d_out[49]
  PIN d_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 0.000 524.770 4.000 ;
    END
  END d_out[4]
  PIN d_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.330 0.000 687.610 4.000 ;
    END
  END d_out[50]
  PIN d_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.010 0.000 691.290 4.000 ;
    END
  END d_out[51]
  PIN d_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 0.000 694.510 4.000 ;
    END
  END d_out[52]
  PIN d_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.910 0.000 698.190 4.000 ;
    END
  END d_out[53]
  PIN d_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.590 0.000 701.870 4.000 ;
    END
  END d_out[54]
  PIN d_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 4.000 ;
    END
  END d_out[55]
  PIN d_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 0.000 708.770 4.000 ;
    END
  END d_out[56]
  PIN d_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 0.000 712.450 4.000 ;
    END
  END d_out[57]
  PIN d_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 0.000 716.130 4.000 ;
    END
  END d_out[58]
  PIN d_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.070 0.000 719.350 4.000 ;
    END
  END d_out[59]
  PIN d_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END d_out[5]
  PIN d_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.750 0.000 723.030 4.000 ;
    END
  END d_out[60]
  PIN d_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.430 0.000 726.710 4.000 ;
    END
  END d_out[61]
  PIN d_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END d_out[62]
  PIN d_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.330 0.000 733.610 4.000 ;
    END
  END d_out[63]
  PIN d_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 0.000 737.290 4.000 ;
    END
  END d_out[64]
  PIN d_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.230 0.000 740.510 4.000 ;
    END
  END d_out[65]
  PIN d_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END d_out[66]
  PIN d_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.590 0.000 747.870 4.000 ;
    END
  END d_out[67]
  PIN d_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 0.000 532.130 4.000 ;
    END
  END d_out[6]
  PIN d_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 0.000 535.350 4.000 ;
    END
  END d_out[7]
  PIN d_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 0.000 539.030 4.000 ;
    END
  END d_out[8]
  PIN d_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END d_out[9]
  PIN m_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END m_in[0]
  PIN m_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 381.520 4.000 382.120 ;
    END
  END m_in[100]
  PIN m_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 385.600 4.000 386.200 ;
    END
  END m_in[101]
  PIN m_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END m_in[102]
  PIN m_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END m_in[103]
  PIN m_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 396.480 4.000 397.080 ;
    END
  END m_in[104]
  PIN m_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 400.560 4.000 401.160 ;
    END
  END m_in[105]
  PIN m_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END m_in[106]
  PIN m_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END m_in[107]
  PIN m_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END m_in[108]
  PIN m_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 415.520 4.000 416.120 ;
    END
  END m_in[109]
  PIN m_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END m_in[10]
  PIN m_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END m_in[110]
  PIN m_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END m_in[111]
  PIN m_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 426.400 4.000 427.000 ;
    END
  END m_in[112]
  PIN m_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 430.480 4.000 431.080 ;
    END
  END m_in[113]
  PIN m_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END m_in[114]
  PIN m_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END m_in[115]
  PIN m_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 441.360 4.000 441.960 ;
    END
  END m_in[116]
  PIN m_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END m_in[117]
  PIN m_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END m_in[118]
  PIN m_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END m_in[119]
  PIN m_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END m_in[11]
  PIN m_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 456.320 4.000 456.920 ;
    END
  END m_in[120]
  PIN m_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 4.000 460.320 ;
    END
  END m_in[121]
  PIN m_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END m_in[122]
  PIN m_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.200 4.000 467.800 ;
    END
  END m_in[123]
  PIN m_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.280 4.000 471.880 ;
    END
  END m_in[124]
  PIN m_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END m_in[125]
  PIN m_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END m_in[126]
  PIN m_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.160 4.000 482.760 ;
    END
  END m_in[127]
  PIN m_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END m_in[128]
  PIN m_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END m_in[129]
  PIN m_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END m_in[12]
  PIN m_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END m_in[130]
  PIN m_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.120 4.000 497.720 ;
    END
  END m_in[131]
  PIN m_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END m_in[13]
  PIN m_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END m_in[14]
  PIN m_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END m_in[15]
  PIN m_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END m_in[16]
  PIN m_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END m_in[17]
  PIN m_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END m_in[18]
  PIN m_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END m_in[19]
  PIN m_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END m_in[1]
  PIN m_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END m_in[20]
  PIN m_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END m_in[21]
  PIN m_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END m_in[22]
  PIN m_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 4.000 95.160 ;
    END
  END m_in[23]
  PIN m_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END m_in[24]
  PIN m_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END m_in[25]
  PIN m_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END m_in[26]
  PIN m_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END m_in[27]
  PIN m_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END m_in[28]
  PIN m_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END m_in[29]
  PIN m_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END m_in[2]
  PIN m_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END m_in[30]
  PIN m_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END m_in[31]
  PIN m_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END m_in[32]
  PIN m_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END m_in[33]
  PIN m_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 4.000 135.960 ;
    END
  END m_in[34]
  PIN m_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END m_in[35]
  PIN m_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END m_in[36]
  PIN m_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END m_in[37]
  PIN m_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.320 4.000 150.920 ;
    END
  END m_in[38]
  PIN m_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END m_in[39]
  PIN m_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END m_in[3]
  PIN m_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END m_in[40]
  PIN m_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 4.000 161.800 ;
    END
  END m_in[41]
  PIN m_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END m_in[42]
  PIN m_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END m_in[43]
  PIN m_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END m_in[44]
  PIN m_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.160 4.000 176.760 ;
    END
  END m_in[45]
  PIN m_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END m_in[46]
  PIN m_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END m_in[47]
  PIN m_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END m_in[48]
  PIN m_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END m_in[49]
  PIN m_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END m_in[4]
  PIN m_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.200 4.000 195.800 ;
    END
  END m_in[50]
  PIN m_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END m_in[51]
  PIN m_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END m_in[52]
  PIN m_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END m_in[53]
  PIN m_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.160 4.000 210.760 ;
    END
  END m_in[54]
  PIN m_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END m_in[55]
  PIN m_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END m_in[56]
  PIN m_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END m_in[57]
  PIN m_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END m_in[58]
  PIN m_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END m_in[59]
  PIN m_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END m_in[5]
  PIN m_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END m_in[60]
  PIN m_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END m_in[61]
  PIN m_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END m_in[62]
  PIN m_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END m_in[63]
  PIN m_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END m_in[64]
  PIN m_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.960 4.000 251.560 ;
    END
  END m_in[65]
  PIN m_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END m_in[66]
  PIN m_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END m_in[67]
  PIN m_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END m_in[68]
  PIN m_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.920 4.000 266.520 ;
    END
  END m_in[69]
  PIN m_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END m_in[6]
  PIN m_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END m_in[70]
  PIN m_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END m_in[71]
  PIN m_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END m_in[72]
  PIN m_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 4.000 281.480 ;
    END
  END m_in[73]
  PIN m_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.960 4.000 285.560 ;
    END
  END m_in[74]
  PIN m_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END m_in[75]
  PIN m_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END m_in[76]
  PIN m_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END m_in[77]
  PIN m_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.920 4.000 300.520 ;
    END
  END m_in[78]
  PIN m_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END m_in[79]
  PIN m_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END m_in[7]
  PIN m_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.720 4.000 307.320 ;
    END
  END m_in[80]
  PIN m_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.800 4.000 311.400 ;
    END
  END m_in[81]
  PIN m_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END m_in[82]
  PIN m_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END m_in[83]
  PIN m_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.680 4.000 322.280 ;
    END
  END m_in[84]
  PIN m_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END m_in[85]
  PIN m_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END m_in[86]
  PIN m_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END m_in[87]
  PIN m_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END m_in[88]
  PIN m_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END m_in[89]
  PIN m_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END m_in[8]
  PIN m_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END m_in[90]
  PIN m_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 4.000 348.800 ;
    END
  END m_in[91]
  PIN m_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.600 4.000 352.200 ;
    END
  END m_in[92]
  PIN m_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.680 4.000 356.280 ;
    END
  END m_in[93]
  PIN m_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END m_in[94]
  PIN m_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END m_in[95]
  PIN m_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.560 4.000 367.160 ;
    END
  END m_in[96]
  PIN m_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END m_in[97]
  PIN m_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END m_in[98]
  PIN m_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END m_in[99]
  PIN m_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END m_in[9]
  PIN m_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.200 4.000 501.800 ;
    END
  END m_out[0]
  PIN m_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 538.600 4.000 539.200 ;
    END
  END m_out[10]
  PIN m_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.000 4.000 542.600 ;
    END
  END m_out[11]
  PIN m_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.080 4.000 546.680 ;
    END
  END m_out[12]
  PIN m_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 549.480 4.000 550.080 ;
    END
  END m_out[13]
  PIN m_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 553.560 4.000 554.160 ;
    END
  END m_out[14]
  PIN m_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.960 4.000 557.560 ;
    END
  END m_out[15]
  PIN m_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END m_out[16]
  PIN m_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END m_out[17]
  PIN m_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 568.520 4.000 569.120 ;
    END
  END m_out[18]
  PIN m_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.920 4.000 572.520 ;
    END
  END m_out[19]
  PIN m_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END m_out[1]
  PIN m_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 576.000 4.000 576.600 ;
    END
  END m_out[20]
  PIN m_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 579.400 4.000 580.000 ;
    END
  END m_out[21]
  PIN m_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END m_out[22]
  PIN m_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.880 4.000 587.480 ;
    END
  END m_out[23]
  PIN m_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.960 4.000 591.560 ;
    END
  END m_out[24]
  PIN m_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 594.360 4.000 594.960 ;
    END
  END m_out[25]
  PIN m_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END m_out[26]
  PIN m_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 4.000 602.440 ;
    END
  END m_out[27]
  PIN m_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END m_out[28]
  PIN m_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 609.320 4.000 609.920 ;
    END
  END m_out[29]
  PIN m_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.680 4.000 509.280 ;
    END
  END m_out[2]
  PIN m_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.720 4.000 613.320 ;
    END
  END m_out[30]
  PIN m_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.800 4.000 617.400 ;
    END
  END m_out[31]
  PIN m_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.200 4.000 620.800 ;
    END
  END m_out[32]
  PIN m_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END m_out[33]
  PIN m_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.680 4.000 628.280 ;
    END
  END m_out[34]
  PIN m_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.760 4.000 632.360 ;
    END
  END m_out[35]
  PIN m_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.160 4.000 635.760 ;
    END
  END m_out[36]
  PIN m_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END m_out[37]
  PIN m_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END m_out[38]
  PIN m_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.720 4.000 647.320 ;
    END
  END m_out[39]
  PIN m_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.080 4.000 512.680 ;
    END
  END m_out[3]
  PIN m_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.120 4.000 650.720 ;
    END
  END m_out[40]
  PIN m_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.200 4.000 654.800 ;
    END
  END m_out[41]
  PIN m_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 657.600 4.000 658.200 ;
    END
  END m_out[42]
  PIN m_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.680 4.000 662.280 ;
    END
  END m_out[43]
  PIN m_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.080 4.000 665.680 ;
    END
  END m_out[44]
  PIN m_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.160 4.000 669.760 ;
    END
  END m_out[45]
  PIN m_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 672.560 4.000 673.160 ;
    END
  END m_out[46]
  PIN m_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 4.000 677.240 ;
    END
  END m_out[47]
  PIN m_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END m_out[48]
  PIN m_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END m_out[49]
  PIN m_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.160 4.000 516.760 ;
    END
  END m_out[4]
  PIN m_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 687.520 4.000 688.120 ;
    END
  END m_out[50]
  PIN m_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 691.600 4.000 692.200 ;
    END
  END m_out[51]
  PIN m_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.000 4.000 695.600 ;
    END
  END m_out[52]
  PIN m_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.080 4.000 699.680 ;
    END
  END m_out[53]
  PIN m_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 702.480 4.000 703.080 ;
    END
  END m_out[54]
  PIN m_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 706.560 4.000 707.160 ;
    END
  END m_out[55]
  PIN m_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 709.960 4.000 710.560 ;
    END
  END m_out[56]
  PIN m_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END m_out[57]
  PIN m_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END m_out[58]
  PIN m_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 721.520 4.000 722.120 ;
    END
  END m_out[59]
  PIN m_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END m_out[5]
  PIN m_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.920 4.000 725.520 ;
    END
  END m_out[60]
  PIN m_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 729.000 4.000 729.600 ;
    END
  END m_out[61]
  PIN m_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 732.400 4.000 733.000 ;
    END
  END m_out[62]
  PIN m_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 736.480 4.000 737.080 ;
    END
  END m_out[63]
  PIN m_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 739.880 4.000 740.480 ;
    END
  END m_out[64]
  PIN m_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.960 4.000 744.560 ;
    END
  END m_out[65]
  PIN m_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 747.360 4.000 747.960 ;
    END
  END m_out[66]
  PIN m_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END m_out[6]
  PIN m_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END m_out[7]
  PIN m_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.120 4.000 531.720 ;
    END
  END m_out[8]
  PIN m_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 534.520 4.000 535.120 ;
    END
  END m_out[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END rst
  PIN stall_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END stall_out
  PIN wishbone_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 746.000 2.210 750.000 ;
    END
  END wishbone_in[0]
  PIN wishbone_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 746.000 45.450 750.000 ;
    END
  END wishbone_in[10]
  PIN wishbone_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 746.000 49.590 750.000 ;
    END
  END wishbone_in[11]
  PIN wishbone_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 746.000 54.190 750.000 ;
    END
  END wishbone_in[12]
  PIN wishbone_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 746.000 58.330 750.000 ;
    END
  END wishbone_in[13]
  PIN wishbone_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 746.000 62.470 750.000 ;
    END
  END wishbone_in[14]
  PIN wishbone_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 746.000 67.070 750.000 ;
    END
  END wishbone_in[15]
  PIN wishbone_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 746.000 71.210 750.000 ;
    END
  END wishbone_in[16]
  PIN wishbone_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 746.000 75.810 750.000 ;
    END
  END wishbone_in[17]
  PIN wishbone_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 746.000 79.950 750.000 ;
    END
  END wishbone_in[18]
  PIN wishbone_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 746.000 84.550 750.000 ;
    END
  END wishbone_in[19]
  PIN wishbone_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 746.000 6.350 750.000 ;
    END
  END wishbone_in[1]
  PIN wishbone_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 746.000 88.690 750.000 ;
    END
  END wishbone_in[20]
  PIN wishbone_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 746.000 92.830 750.000 ;
    END
  END wishbone_in[21]
  PIN wishbone_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 746.000 97.430 750.000 ;
    END
  END wishbone_in[22]
  PIN wishbone_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 746.000 101.570 750.000 ;
    END
  END wishbone_in[23]
  PIN wishbone_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 746.000 106.170 750.000 ;
    END
  END wishbone_in[24]
  PIN wishbone_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 746.000 110.310 750.000 ;
    END
  END wishbone_in[25]
  PIN wishbone_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 746.000 114.450 750.000 ;
    END
  END wishbone_in[26]
  PIN wishbone_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 746.000 119.050 750.000 ;
    END
  END wishbone_in[27]
  PIN wishbone_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 746.000 123.190 750.000 ;
    END
  END wishbone_in[28]
  PIN wishbone_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 746.000 127.790 750.000 ;
    END
  END wishbone_in[29]
  PIN wishbone_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 746.000 10.490 750.000 ;
    END
  END wishbone_in[2]
  PIN wishbone_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 746.000 131.930 750.000 ;
    END
  END wishbone_in[30]
  PIN wishbone_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 746.000 136.530 750.000 ;
    END
  END wishbone_in[31]
  PIN wishbone_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 746.000 140.670 750.000 ;
    END
  END wishbone_in[32]
  PIN wishbone_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 746.000 144.810 750.000 ;
    END
  END wishbone_in[33]
  PIN wishbone_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 746.000 149.410 750.000 ;
    END
  END wishbone_in[34]
  PIN wishbone_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 746.000 153.550 750.000 ;
    END
  END wishbone_in[35]
  PIN wishbone_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 746.000 158.150 750.000 ;
    END
  END wishbone_in[36]
  PIN wishbone_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 746.000 162.290 750.000 ;
    END
  END wishbone_in[37]
  PIN wishbone_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 746.000 166.890 750.000 ;
    END
  END wishbone_in[38]
  PIN wishbone_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 746.000 171.030 750.000 ;
    END
  END wishbone_in[39]
  PIN wishbone_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 746.000 15.090 750.000 ;
    END
  END wishbone_in[3]
  PIN wishbone_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 746.000 175.170 750.000 ;
    END
  END wishbone_in[40]
  PIN wishbone_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 746.000 179.770 750.000 ;
    END
  END wishbone_in[41]
  PIN wishbone_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 746.000 183.910 750.000 ;
    END
  END wishbone_in[42]
  PIN wishbone_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 746.000 188.510 750.000 ;
    END
  END wishbone_in[43]
  PIN wishbone_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 746.000 192.650 750.000 ;
    END
  END wishbone_in[44]
  PIN wishbone_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 746.000 196.790 750.000 ;
    END
  END wishbone_in[45]
  PIN wishbone_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 746.000 201.390 750.000 ;
    END
  END wishbone_in[46]
  PIN wishbone_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 746.000 205.530 750.000 ;
    END
  END wishbone_in[47]
  PIN wishbone_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 746.000 210.130 750.000 ;
    END
  END wishbone_in[48]
  PIN wishbone_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 746.000 214.270 750.000 ;
    END
  END wishbone_in[49]
  PIN wishbone_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 746.000 19.230 750.000 ;
    END
  END wishbone_in[4]
  PIN wishbone_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 746.000 218.870 750.000 ;
    END
  END wishbone_in[50]
  PIN wishbone_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 746.000 223.010 750.000 ;
    END
  END wishbone_in[51]
  PIN wishbone_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 746.000 227.150 750.000 ;
    END
  END wishbone_in[52]
  PIN wishbone_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 746.000 231.750 750.000 ;
    END
  END wishbone_in[53]
  PIN wishbone_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 746.000 235.890 750.000 ;
    END
  END wishbone_in[54]
  PIN wishbone_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 746.000 240.490 750.000 ;
    END
  END wishbone_in[55]
  PIN wishbone_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 746.000 244.630 750.000 ;
    END
  END wishbone_in[56]
  PIN wishbone_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 746.000 249.230 750.000 ;
    END
  END wishbone_in[57]
  PIN wishbone_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 746.000 253.370 750.000 ;
    END
  END wishbone_in[58]
  PIN wishbone_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 746.000 257.510 750.000 ;
    END
  END wishbone_in[59]
  PIN wishbone_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 746.000 23.830 750.000 ;
    END
  END wishbone_in[5]
  PIN wishbone_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 746.000 262.110 750.000 ;
    END
  END wishbone_in[60]
  PIN wishbone_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 746.000 266.250 750.000 ;
    END
  END wishbone_in[61]
  PIN wishbone_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 746.000 270.850 750.000 ;
    END
  END wishbone_in[62]
  PIN wishbone_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 746.000 274.990 750.000 ;
    END
  END wishbone_in[63]
  PIN wishbone_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 746.000 279.590 750.000 ;
    END
  END wishbone_in[64]
  PIN wishbone_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 746.000 283.730 750.000 ;
    END
  END wishbone_in[65]
  PIN wishbone_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 746.000 27.970 750.000 ;
    END
  END wishbone_in[6]
  PIN wishbone_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 746.000 32.110 750.000 ;
    END
  END wishbone_in[7]
  PIN wishbone_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 746.000 36.710 750.000 ;
    END
  END wishbone_in[8]
  PIN wishbone_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 746.000 40.850 750.000 ;
    END
  END wishbone_in[9]
  PIN wishbone_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 746.000 287.870 750.000 ;
    END
  END wishbone_out[0]
  PIN wishbone_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 746.000 721.650 750.000 ;
    END
  END wishbone_out[100]
  PIN wishbone_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.510 746.000 725.790 750.000 ;
    END
  END wishbone_out[101]
  PIN wishbone_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 746.000 729.930 750.000 ;
    END
  END wishbone_out[102]
  PIN wishbone_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 746.000 734.530 750.000 ;
    END
  END wishbone_out[103]
  PIN wishbone_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.390 746.000 738.670 750.000 ;
    END
  END wishbone_out[104]
  PIN wishbone_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.990 746.000 743.270 750.000 ;
    END
  END wishbone_out[105]
  PIN wishbone_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 746.000 747.410 750.000 ;
    END
  END wishbone_out[106]
  PIN wishbone_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 746.000 331.570 750.000 ;
    END
  END wishbone_out[10]
  PIN wishbone_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 746.000 335.710 750.000 ;
    END
  END wishbone_out[11]
  PIN wishbone_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 746.000 339.850 750.000 ;
    END
  END wishbone_out[12]
  PIN wishbone_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 746.000 344.450 750.000 ;
    END
  END wishbone_out[13]
  PIN wishbone_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 746.000 348.590 750.000 ;
    END
  END wishbone_out[14]
  PIN wishbone_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 746.000 353.190 750.000 ;
    END
  END wishbone_out[15]
  PIN wishbone_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 746.000 357.330 750.000 ;
    END
  END wishbone_out[16]
  PIN wishbone_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 746.000 361.930 750.000 ;
    END
  END wishbone_out[17]
  PIN wishbone_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 746.000 366.070 750.000 ;
    END
  END wishbone_out[18]
  PIN wishbone_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 746.000 370.210 750.000 ;
    END
  END wishbone_out[19]
  PIN wishbone_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 746.000 292.470 750.000 ;
    END
  END wishbone_out[1]
  PIN wishbone_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 746.000 374.810 750.000 ;
    END
  END wishbone_out[20]
  PIN wishbone_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 746.000 378.950 750.000 ;
    END
  END wishbone_out[21]
  PIN wishbone_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 746.000 383.550 750.000 ;
    END
  END wishbone_out[22]
  PIN wishbone_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.410 746.000 387.690 750.000 ;
    END
  END wishbone_out[23]
  PIN wishbone_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 746.000 391.830 750.000 ;
    END
  END wishbone_out[24]
  PIN wishbone_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 746.000 396.430 750.000 ;
    END
  END wishbone_out[25]
  PIN wishbone_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 746.000 400.570 750.000 ;
    END
  END wishbone_out[26]
  PIN wishbone_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 746.000 405.170 750.000 ;
    END
  END wishbone_out[27]
  PIN wishbone_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 746.000 409.310 750.000 ;
    END
  END wishbone_out[28]
  PIN wishbone_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 746.000 413.910 750.000 ;
    END
  END wishbone_out[29]
  PIN wishbone_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 746.000 296.610 750.000 ;
    END
  END wishbone_out[2]
  PIN wishbone_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 746.000 418.050 750.000 ;
    END
  END wishbone_out[30]
  PIN wishbone_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 746.000 422.190 750.000 ;
    END
  END wishbone_out[31]
  PIN wishbone_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 746.000 426.790 750.000 ;
    END
  END wishbone_out[32]
  PIN wishbone_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 746.000 430.930 750.000 ;
    END
  END wishbone_out[33]
  PIN wishbone_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 746.000 435.530 750.000 ;
    END
  END wishbone_out[34]
  PIN wishbone_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 746.000 439.670 750.000 ;
    END
  END wishbone_out[35]
  PIN wishbone_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 746.000 444.270 750.000 ;
    END
  END wishbone_out[36]
  PIN wishbone_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.130 746.000 448.410 750.000 ;
    END
  END wishbone_out[37]
  PIN wishbone_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 746.000 452.550 750.000 ;
    END
  END wishbone_out[38]
  PIN wishbone_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 746.000 457.150 750.000 ;
    END
  END wishbone_out[39]
  PIN wishbone_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 746.000 301.210 750.000 ;
    END
  END wishbone_out[3]
  PIN wishbone_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 746.000 461.290 750.000 ;
    END
  END wishbone_out[40]
  PIN wishbone_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 746.000 465.890 750.000 ;
    END
  END wishbone_out[41]
  PIN wishbone_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 746.000 470.030 750.000 ;
    END
  END wishbone_out[42]
  PIN wishbone_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 746.000 474.170 750.000 ;
    END
  END wishbone_out[43]
  PIN wishbone_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 746.000 478.770 750.000 ;
    END
  END wishbone_out[44]
  PIN wishbone_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 746.000 482.910 750.000 ;
    END
  END wishbone_out[45]
  PIN wishbone_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 746.000 487.510 750.000 ;
    END
  END wishbone_out[46]
  PIN wishbone_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 746.000 491.650 750.000 ;
    END
  END wishbone_out[47]
  PIN wishbone_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 746.000 496.250 750.000 ;
    END
  END wishbone_out[48]
  PIN wishbone_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.110 746.000 500.390 750.000 ;
    END
  END wishbone_out[49]
  PIN wishbone_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 746.000 305.350 750.000 ;
    END
  END wishbone_out[4]
  PIN wishbone_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 746.000 504.530 750.000 ;
    END
  END wishbone_out[50]
  PIN wishbone_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 746.000 509.130 750.000 ;
    END
  END wishbone_out[51]
  PIN wishbone_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 746.000 513.270 750.000 ;
    END
  END wishbone_out[52]
  PIN wishbone_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 746.000 517.870 750.000 ;
    END
  END wishbone_out[53]
  PIN wishbone_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 746.000 522.010 750.000 ;
    END
  END wishbone_out[54]
  PIN wishbone_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 746.000 526.610 750.000 ;
    END
  END wishbone_out[55]
  PIN wishbone_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 746.000 530.750 750.000 ;
    END
  END wishbone_out[56]
  PIN wishbone_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 746.000 534.890 750.000 ;
    END
  END wishbone_out[57]
  PIN wishbone_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 746.000 539.490 750.000 ;
    END
  END wishbone_out[58]
  PIN wishbone_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 746.000 543.630 750.000 ;
    END
  END wishbone_out[59]
  PIN wishbone_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 746.000 309.490 750.000 ;
    END
  END wishbone_out[5]
  PIN wishbone_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 746.000 548.230 750.000 ;
    END
  END wishbone_out[60]
  PIN wishbone_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 746.000 552.370 750.000 ;
    END
  END wishbone_out[61]
  PIN wishbone_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 746.000 556.970 750.000 ;
    END
  END wishbone_out[62]
  PIN wishbone_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 746.000 561.110 750.000 ;
    END
  END wishbone_out[63]
  PIN wishbone_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 746.000 565.250 750.000 ;
    END
  END wishbone_out[64]
  PIN wishbone_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 746.000 569.850 750.000 ;
    END
  END wishbone_out[65]
  PIN wishbone_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.710 746.000 573.990 750.000 ;
    END
  END wishbone_out[66]
  PIN wishbone_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 746.000 578.590 750.000 ;
    END
  END wishbone_out[67]
  PIN wishbone_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 746.000 582.730 750.000 ;
    END
  END wishbone_out[68]
  PIN wishbone_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 746.000 586.870 750.000 ;
    END
  END wishbone_out[69]
  PIN wishbone_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 746.000 314.090 750.000 ;
    END
  END wishbone_out[6]
  PIN wishbone_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 746.000 591.470 750.000 ;
    END
  END wishbone_out[70]
  PIN wishbone_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 746.000 595.610 750.000 ;
    END
  END wishbone_out[71]
  PIN wishbone_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 746.000 600.210 750.000 ;
    END
  END wishbone_out[72]
  PIN wishbone_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 746.000 604.350 750.000 ;
    END
  END wishbone_out[73]
  PIN wishbone_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 746.000 608.950 750.000 ;
    END
  END wishbone_out[74]
  PIN wishbone_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 746.000 613.090 750.000 ;
    END
  END wishbone_out[75]
  PIN wishbone_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.950 746.000 617.230 750.000 ;
    END
  END wishbone_out[76]
  PIN wishbone_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 746.000 621.830 750.000 ;
    END
  END wishbone_out[77]
  PIN wishbone_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 746.000 625.970 750.000 ;
    END
  END wishbone_out[78]
  PIN wishbone_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 746.000 630.570 750.000 ;
    END
  END wishbone_out[79]
  PIN wishbone_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 746.000 318.230 750.000 ;
    END
  END wishbone_out[7]
  PIN wishbone_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 746.000 634.710 750.000 ;
    END
  END wishbone_out[80]
  PIN wishbone_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 746.000 639.310 750.000 ;
    END
  END wishbone_out[81]
  PIN wishbone_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 746.000 643.450 750.000 ;
    END
  END wishbone_out[82]
  PIN wishbone_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 746.000 647.590 750.000 ;
    END
  END wishbone_out[83]
  PIN wishbone_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.910 746.000 652.190 750.000 ;
    END
  END wishbone_out[84]
  PIN wishbone_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.050 746.000 656.330 750.000 ;
    END
  END wishbone_out[85]
  PIN wishbone_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 746.000 660.930 750.000 ;
    END
  END wishbone_out[86]
  PIN wishbone_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.790 746.000 665.070 750.000 ;
    END
  END wishbone_out[87]
  PIN wishbone_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 746.000 669.210 750.000 ;
    END
  END wishbone_out[88]
  PIN wishbone_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 746.000 673.810 750.000 ;
    END
  END wishbone_out[89]
  PIN wishbone_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 746.000 322.830 750.000 ;
    END
  END wishbone_out[8]
  PIN wishbone_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.670 746.000 677.950 750.000 ;
    END
  END wishbone_out[90]
  PIN wishbone_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.270 746.000 682.550 750.000 ;
    END
  END wishbone_out[91]
  PIN wishbone_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 746.000 686.690 750.000 ;
    END
  END wishbone_out[92]
  PIN wishbone_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.010 746.000 691.290 750.000 ;
    END
  END wishbone_out[93]
  PIN wishbone_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.150 746.000 695.430 750.000 ;
    END
  END wishbone_out[94]
  PIN wishbone_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 746.000 699.570 750.000 ;
    END
  END wishbone_out[95]
  PIN wishbone_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 746.000 704.170 750.000 ;
    END
  END wishbone_out[96]
  PIN wishbone_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.030 746.000 708.310 750.000 ;
    END
  END wishbone_out[97]
  PIN wishbone_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 746.000 712.910 750.000 ;
    END
  END wishbone_out[98]
  PIN wishbone_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.770 746.000 717.050 750.000 ;
    END
  END wishbone_out[99]
  PIN wishbone_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 746.000 326.970 750.000 ;
    END
  END wishbone_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 737.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 737.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 737.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 737.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 737.360 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 737.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 737.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 737.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 737.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 737.360 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 638.740 10.880 640.340 737.120 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 485.140 10.880 486.740 737.120 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 737.120 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 737.120 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 737.120 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 715.540 10.880 717.140 737.120 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 561.940 10.880 563.540 737.120 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 408.340 10.880 409.940 737.120 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 737.120 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 737.120 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 642.040 10.880 643.640 737.120 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 488.440 10.880 490.040 737.120 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.840 10.880 336.440 737.120 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 737.120 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 737.120 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 718.840 10.880 720.440 737.120 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 565.240 10.880 566.840 737.120 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 411.640 10.880 413.240 737.120 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 737.120 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 737.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 645.340 10.880 646.940 737.120 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 491.740 10.880 493.340 737.120 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 338.140 10.880 339.740 737.120 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 737.120 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 737.120 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 722.140 10.880 723.740 737.120 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 568.540 10.880 570.140 737.120 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 414.940 10.880 416.540 737.120 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 737.120 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 737.120 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 7.225 744.280 742.135 ;
      LAYER met1 ;
        RECT 1.450 6.500 747.890 750.000 ;
      LAYER met2 ;
        RECT 1.480 745.720 1.650 750.030 ;
        RECT 2.490 745.720 5.790 750.030 ;
        RECT 6.630 745.720 9.930 750.030 ;
        RECT 10.770 745.720 14.530 750.030 ;
        RECT 15.370 745.720 18.670 750.030 ;
        RECT 19.510 745.720 23.270 750.030 ;
        RECT 24.110 745.720 27.410 750.030 ;
        RECT 28.250 745.720 31.550 750.030 ;
        RECT 32.390 745.720 36.150 750.030 ;
        RECT 36.990 745.720 40.290 750.030 ;
        RECT 41.130 745.720 44.890 750.030 ;
        RECT 45.730 745.720 49.030 750.030 ;
        RECT 49.870 745.720 53.630 750.030 ;
        RECT 54.470 745.720 57.770 750.030 ;
        RECT 58.610 745.720 61.910 750.030 ;
        RECT 62.750 745.720 66.510 750.030 ;
        RECT 67.350 745.720 70.650 750.030 ;
        RECT 71.490 745.720 75.250 750.030 ;
        RECT 76.090 745.720 79.390 750.030 ;
        RECT 80.230 745.720 83.990 750.030 ;
        RECT 84.830 745.720 88.130 750.030 ;
        RECT 88.970 745.720 92.270 750.030 ;
        RECT 93.110 745.720 96.870 750.030 ;
        RECT 97.710 745.720 101.010 750.030 ;
        RECT 101.850 745.720 105.610 750.030 ;
        RECT 106.450 745.720 109.750 750.030 ;
        RECT 110.590 745.720 113.890 750.030 ;
        RECT 114.730 745.720 118.490 750.030 ;
        RECT 119.330 745.720 122.630 750.030 ;
        RECT 123.470 745.720 127.230 750.030 ;
        RECT 128.070 745.720 131.370 750.030 ;
        RECT 132.210 745.720 135.970 750.030 ;
        RECT 136.810 745.720 140.110 750.030 ;
        RECT 140.950 745.720 144.250 750.030 ;
        RECT 145.090 745.720 148.850 750.030 ;
        RECT 149.690 745.720 152.990 750.030 ;
        RECT 153.830 745.720 157.590 750.030 ;
        RECT 158.430 745.720 161.730 750.030 ;
        RECT 162.570 745.720 166.330 750.030 ;
        RECT 167.170 745.720 170.470 750.030 ;
        RECT 171.310 745.720 174.610 750.030 ;
        RECT 175.450 745.720 179.210 750.030 ;
        RECT 180.050 745.720 183.350 750.030 ;
        RECT 184.190 745.720 187.950 750.030 ;
        RECT 188.790 745.720 192.090 750.030 ;
        RECT 192.930 745.720 196.230 750.030 ;
        RECT 197.070 745.720 200.830 750.030 ;
        RECT 201.670 745.720 204.970 750.030 ;
        RECT 205.810 745.720 209.570 750.030 ;
        RECT 210.410 745.720 213.710 750.030 ;
        RECT 214.550 745.720 218.310 750.030 ;
        RECT 219.150 745.720 222.450 750.030 ;
        RECT 223.290 745.720 226.590 750.030 ;
        RECT 227.430 745.720 231.190 750.030 ;
        RECT 232.030 745.720 235.330 750.030 ;
        RECT 236.170 745.720 239.930 750.030 ;
        RECT 240.770 745.720 244.070 750.030 ;
        RECT 244.910 745.720 248.670 750.030 ;
        RECT 249.510 745.720 252.810 750.030 ;
        RECT 253.650 745.720 256.950 750.030 ;
        RECT 257.790 745.720 261.550 750.030 ;
        RECT 262.390 745.720 265.690 750.030 ;
        RECT 266.530 745.720 270.290 750.030 ;
        RECT 271.130 745.720 274.430 750.030 ;
        RECT 275.270 745.720 279.030 750.030 ;
        RECT 279.870 745.720 283.170 750.030 ;
        RECT 284.010 745.720 287.310 750.030 ;
        RECT 288.150 745.720 291.910 750.030 ;
        RECT 292.750 745.720 296.050 750.030 ;
        RECT 296.890 745.720 300.650 750.030 ;
        RECT 301.490 745.720 304.790 750.030 ;
        RECT 305.630 745.720 308.930 750.030 ;
        RECT 309.770 745.720 313.530 750.030 ;
        RECT 314.370 745.720 317.670 750.030 ;
        RECT 318.510 745.720 322.270 750.030 ;
        RECT 323.110 745.720 326.410 750.030 ;
        RECT 327.250 745.720 331.010 750.030 ;
        RECT 331.850 745.720 335.150 750.030 ;
        RECT 335.990 745.720 339.290 750.030 ;
        RECT 340.130 745.720 343.890 750.030 ;
        RECT 344.730 745.720 348.030 750.030 ;
        RECT 348.870 745.720 352.630 750.030 ;
        RECT 353.470 745.720 356.770 750.030 ;
        RECT 357.610 745.720 361.370 750.030 ;
        RECT 362.210 745.720 365.510 750.030 ;
        RECT 366.350 745.720 369.650 750.030 ;
        RECT 370.490 745.720 374.250 750.030 ;
        RECT 375.090 745.720 378.390 750.030 ;
        RECT 379.230 745.720 382.990 750.030 ;
        RECT 383.830 745.720 387.130 750.030 ;
        RECT 387.970 745.720 391.270 750.030 ;
        RECT 392.110 745.720 395.870 750.030 ;
        RECT 396.710 745.720 400.010 750.030 ;
        RECT 400.850 745.720 404.610 750.030 ;
        RECT 405.450 745.720 408.750 750.030 ;
        RECT 409.590 745.720 413.350 750.030 ;
        RECT 414.190 745.720 417.490 750.030 ;
        RECT 418.330 745.720 421.630 750.030 ;
        RECT 422.470 745.720 426.230 750.030 ;
        RECT 427.070 745.720 430.370 750.030 ;
        RECT 431.210 745.720 434.970 750.030 ;
        RECT 435.810 745.720 439.110 750.030 ;
        RECT 439.950 745.720 443.710 750.030 ;
        RECT 444.550 745.720 447.850 750.030 ;
        RECT 448.690 745.720 451.990 750.030 ;
        RECT 452.830 745.720 456.590 750.030 ;
        RECT 457.430 745.720 460.730 750.030 ;
        RECT 461.570 745.720 465.330 750.030 ;
        RECT 466.170 745.720 469.470 750.030 ;
        RECT 470.310 745.720 473.610 750.030 ;
        RECT 474.450 745.720 478.210 750.030 ;
        RECT 479.050 745.720 482.350 750.030 ;
        RECT 483.190 745.720 486.950 750.030 ;
        RECT 487.790 745.720 491.090 750.030 ;
        RECT 491.930 745.720 495.690 750.030 ;
        RECT 496.530 745.720 499.830 750.030 ;
        RECT 500.670 745.720 503.970 750.030 ;
        RECT 504.810 745.720 508.570 750.030 ;
        RECT 509.410 745.720 512.710 750.030 ;
        RECT 513.550 745.720 517.310 750.030 ;
        RECT 518.150 745.720 521.450 750.030 ;
        RECT 522.290 745.720 526.050 750.030 ;
        RECT 526.890 745.720 530.190 750.030 ;
        RECT 531.030 745.720 534.330 750.030 ;
        RECT 535.170 745.720 538.930 750.030 ;
        RECT 539.770 745.720 543.070 750.030 ;
        RECT 543.910 745.720 547.670 750.030 ;
        RECT 548.510 745.720 551.810 750.030 ;
        RECT 552.650 745.720 556.410 750.030 ;
        RECT 557.250 745.720 560.550 750.030 ;
        RECT 561.390 745.720 564.690 750.030 ;
        RECT 565.530 745.720 569.290 750.030 ;
        RECT 570.130 745.720 573.430 750.030 ;
        RECT 574.270 745.720 578.030 750.030 ;
        RECT 578.870 745.720 582.170 750.030 ;
        RECT 583.010 745.720 586.310 750.030 ;
        RECT 587.150 745.720 590.910 750.030 ;
        RECT 591.750 745.720 595.050 750.030 ;
        RECT 595.890 745.720 599.650 750.030 ;
        RECT 600.490 745.720 603.790 750.030 ;
        RECT 604.630 745.720 608.390 750.030 ;
        RECT 609.230 745.720 612.530 750.030 ;
        RECT 613.370 745.720 616.670 750.030 ;
        RECT 617.510 745.720 621.270 750.030 ;
        RECT 622.110 745.720 625.410 750.030 ;
        RECT 626.250 745.720 630.010 750.030 ;
        RECT 630.850 745.720 634.150 750.030 ;
        RECT 634.990 745.720 638.750 750.030 ;
        RECT 639.590 745.720 642.890 750.030 ;
        RECT 643.730 745.720 647.030 750.030 ;
        RECT 647.870 745.720 651.630 750.030 ;
        RECT 652.470 745.720 655.770 750.030 ;
        RECT 656.610 745.720 660.370 750.030 ;
        RECT 661.210 745.720 664.510 750.030 ;
        RECT 665.350 745.720 668.650 750.030 ;
        RECT 669.490 745.720 673.250 750.030 ;
        RECT 674.090 745.720 677.390 750.030 ;
        RECT 678.230 745.720 681.990 750.030 ;
        RECT 682.830 745.720 686.130 750.030 ;
        RECT 686.970 745.720 690.730 750.030 ;
        RECT 691.570 745.720 694.870 750.030 ;
        RECT 695.710 745.720 699.010 750.030 ;
        RECT 699.850 745.720 703.610 750.030 ;
        RECT 704.450 745.720 707.750 750.030 ;
        RECT 708.590 745.720 712.350 750.030 ;
        RECT 713.190 745.720 716.490 750.030 ;
        RECT 717.330 745.720 721.090 750.030 ;
        RECT 721.930 745.720 725.230 750.030 ;
        RECT 726.070 745.720 729.370 750.030 ;
        RECT 730.210 745.720 733.970 750.030 ;
        RECT 734.810 745.720 738.110 750.030 ;
        RECT 738.950 745.720 742.710 750.030 ;
        RECT 743.550 745.720 746.850 750.030 ;
        RECT 747.690 745.720 747.860 750.030 ;
        RECT 1.480 4.280 747.860 745.720 ;
        RECT 2.030 4.000 4.410 4.280 ;
        RECT 5.250 4.000 8.090 4.280 ;
        RECT 8.930 4.000 11.770 4.280 ;
        RECT 12.610 4.000 14.990 4.280 ;
        RECT 15.830 4.000 18.670 4.280 ;
        RECT 19.510 4.000 22.350 4.280 ;
        RECT 23.190 4.000 25.570 4.280 ;
        RECT 26.410 4.000 29.250 4.280 ;
        RECT 30.090 4.000 32.930 4.280 ;
        RECT 33.770 4.000 36.150 4.280 ;
        RECT 36.990 4.000 39.830 4.280 ;
        RECT 40.670 4.000 43.510 4.280 ;
        RECT 44.350 4.000 46.730 4.280 ;
        RECT 47.570 4.000 50.410 4.280 ;
        RECT 51.250 4.000 54.090 4.280 ;
        RECT 54.930 4.000 57.770 4.280 ;
        RECT 58.610 4.000 60.990 4.280 ;
        RECT 61.830 4.000 64.670 4.280 ;
        RECT 65.510 4.000 68.350 4.280 ;
        RECT 69.190 4.000 71.570 4.280 ;
        RECT 72.410 4.000 75.250 4.280 ;
        RECT 76.090 4.000 78.930 4.280 ;
        RECT 79.770 4.000 82.150 4.280 ;
        RECT 82.990 4.000 85.830 4.280 ;
        RECT 86.670 4.000 89.510 4.280 ;
        RECT 90.350 4.000 92.730 4.280 ;
        RECT 93.570 4.000 96.410 4.280 ;
        RECT 97.250 4.000 100.090 4.280 ;
        RECT 100.930 4.000 103.310 4.280 ;
        RECT 104.150 4.000 106.990 4.280 ;
        RECT 107.830 4.000 110.670 4.280 ;
        RECT 111.510 4.000 114.350 4.280 ;
        RECT 115.190 4.000 117.570 4.280 ;
        RECT 118.410 4.000 121.250 4.280 ;
        RECT 122.090 4.000 124.930 4.280 ;
        RECT 125.770 4.000 128.150 4.280 ;
        RECT 128.990 4.000 131.830 4.280 ;
        RECT 132.670 4.000 135.510 4.280 ;
        RECT 136.350 4.000 138.730 4.280 ;
        RECT 139.570 4.000 142.410 4.280 ;
        RECT 143.250 4.000 146.090 4.280 ;
        RECT 146.930 4.000 149.310 4.280 ;
        RECT 150.150 4.000 152.990 4.280 ;
        RECT 153.830 4.000 156.670 4.280 ;
        RECT 157.510 4.000 159.890 4.280 ;
        RECT 160.730 4.000 163.570 4.280 ;
        RECT 164.410 4.000 167.250 4.280 ;
        RECT 168.090 4.000 170.930 4.280 ;
        RECT 171.770 4.000 174.150 4.280 ;
        RECT 174.990 4.000 177.830 4.280 ;
        RECT 178.670 4.000 181.510 4.280 ;
        RECT 182.350 4.000 184.730 4.280 ;
        RECT 185.570 4.000 188.410 4.280 ;
        RECT 189.250 4.000 192.090 4.280 ;
        RECT 192.930 4.000 195.310 4.280 ;
        RECT 196.150 4.000 198.990 4.280 ;
        RECT 199.830 4.000 202.670 4.280 ;
        RECT 203.510 4.000 205.890 4.280 ;
        RECT 206.730 4.000 209.570 4.280 ;
        RECT 210.410 4.000 213.250 4.280 ;
        RECT 214.090 4.000 216.930 4.280 ;
        RECT 217.770 4.000 220.150 4.280 ;
        RECT 220.990 4.000 223.830 4.280 ;
        RECT 224.670 4.000 227.510 4.280 ;
        RECT 228.350 4.000 230.730 4.280 ;
        RECT 231.570 4.000 234.410 4.280 ;
        RECT 235.250 4.000 238.090 4.280 ;
        RECT 238.930 4.000 241.310 4.280 ;
        RECT 242.150 4.000 244.990 4.280 ;
        RECT 245.830 4.000 248.670 4.280 ;
        RECT 249.510 4.000 251.890 4.280 ;
        RECT 252.730 4.000 255.570 4.280 ;
        RECT 256.410 4.000 259.250 4.280 ;
        RECT 260.090 4.000 262.470 4.280 ;
        RECT 263.310 4.000 266.150 4.280 ;
        RECT 266.990 4.000 269.830 4.280 ;
        RECT 270.670 4.000 273.510 4.280 ;
        RECT 274.350 4.000 276.730 4.280 ;
        RECT 277.570 4.000 280.410 4.280 ;
        RECT 281.250 4.000 284.090 4.280 ;
        RECT 284.930 4.000 287.310 4.280 ;
        RECT 288.150 4.000 290.990 4.280 ;
        RECT 291.830 4.000 294.670 4.280 ;
        RECT 295.510 4.000 297.890 4.280 ;
        RECT 298.730 4.000 301.570 4.280 ;
        RECT 302.410 4.000 305.250 4.280 ;
        RECT 306.090 4.000 308.470 4.280 ;
        RECT 309.310 4.000 312.150 4.280 ;
        RECT 312.990 4.000 315.830 4.280 ;
        RECT 316.670 4.000 319.050 4.280 ;
        RECT 319.890 4.000 322.730 4.280 ;
        RECT 323.570 4.000 326.410 4.280 ;
        RECT 327.250 4.000 330.090 4.280 ;
        RECT 330.930 4.000 333.310 4.280 ;
        RECT 334.150 4.000 336.990 4.280 ;
        RECT 337.830 4.000 340.670 4.280 ;
        RECT 341.510 4.000 343.890 4.280 ;
        RECT 344.730 4.000 347.570 4.280 ;
        RECT 348.410 4.000 351.250 4.280 ;
        RECT 352.090 4.000 354.470 4.280 ;
        RECT 355.310 4.000 358.150 4.280 ;
        RECT 358.990 4.000 361.830 4.280 ;
        RECT 362.670 4.000 365.050 4.280 ;
        RECT 365.890 4.000 368.730 4.280 ;
        RECT 369.570 4.000 372.410 4.280 ;
        RECT 373.250 4.000 376.090 4.280 ;
        RECT 376.930 4.000 379.310 4.280 ;
        RECT 380.150 4.000 382.990 4.280 ;
        RECT 383.830 4.000 386.670 4.280 ;
        RECT 387.510 4.000 389.890 4.280 ;
        RECT 390.730 4.000 393.570 4.280 ;
        RECT 394.410 4.000 397.250 4.280 ;
        RECT 398.090 4.000 400.470 4.280 ;
        RECT 401.310 4.000 404.150 4.280 ;
        RECT 404.990 4.000 407.830 4.280 ;
        RECT 408.670 4.000 411.050 4.280 ;
        RECT 411.890 4.000 414.730 4.280 ;
        RECT 415.570 4.000 418.410 4.280 ;
        RECT 419.250 4.000 421.630 4.280 ;
        RECT 422.470 4.000 425.310 4.280 ;
        RECT 426.150 4.000 428.990 4.280 ;
        RECT 429.830 4.000 432.670 4.280 ;
        RECT 433.510 4.000 435.890 4.280 ;
        RECT 436.730 4.000 439.570 4.280 ;
        RECT 440.410 4.000 443.250 4.280 ;
        RECT 444.090 4.000 446.470 4.280 ;
        RECT 447.310 4.000 450.150 4.280 ;
        RECT 450.990 4.000 453.830 4.280 ;
        RECT 454.670 4.000 457.050 4.280 ;
        RECT 457.890 4.000 460.730 4.280 ;
        RECT 461.570 4.000 464.410 4.280 ;
        RECT 465.250 4.000 467.630 4.280 ;
        RECT 468.470 4.000 471.310 4.280 ;
        RECT 472.150 4.000 474.990 4.280 ;
        RECT 475.830 4.000 478.210 4.280 ;
        RECT 479.050 4.000 481.890 4.280 ;
        RECT 482.730 4.000 485.570 4.280 ;
        RECT 486.410 4.000 489.250 4.280 ;
        RECT 490.090 4.000 492.470 4.280 ;
        RECT 493.310 4.000 496.150 4.280 ;
        RECT 496.990 4.000 499.830 4.280 ;
        RECT 500.670 4.000 503.050 4.280 ;
        RECT 503.890 4.000 506.730 4.280 ;
        RECT 507.570 4.000 510.410 4.280 ;
        RECT 511.250 4.000 513.630 4.280 ;
        RECT 514.470 4.000 517.310 4.280 ;
        RECT 518.150 4.000 520.990 4.280 ;
        RECT 521.830 4.000 524.210 4.280 ;
        RECT 525.050 4.000 527.890 4.280 ;
        RECT 528.730 4.000 531.570 4.280 ;
        RECT 532.410 4.000 534.790 4.280 ;
        RECT 535.630 4.000 538.470 4.280 ;
        RECT 539.310 4.000 542.150 4.280 ;
        RECT 542.990 4.000 545.830 4.280 ;
        RECT 546.670 4.000 549.050 4.280 ;
        RECT 549.890 4.000 552.730 4.280 ;
        RECT 553.570 4.000 556.410 4.280 ;
        RECT 557.250 4.000 559.630 4.280 ;
        RECT 560.470 4.000 563.310 4.280 ;
        RECT 564.150 4.000 566.990 4.280 ;
        RECT 567.830 4.000 570.210 4.280 ;
        RECT 571.050 4.000 573.890 4.280 ;
        RECT 574.730 4.000 577.570 4.280 ;
        RECT 578.410 4.000 580.790 4.280 ;
        RECT 581.630 4.000 584.470 4.280 ;
        RECT 585.310 4.000 588.150 4.280 ;
        RECT 588.990 4.000 591.830 4.280 ;
        RECT 592.670 4.000 595.050 4.280 ;
        RECT 595.890 4.000 598.730 4.280 ;
        RECT 599.570 4.000 602.410 4.280 ;
        RECT 603.250 4.000 605.630 4.280 ;
        RECT 606.470 4.000 609.310 4.280 ;
        RECT 610.150 4.000 612.990 4.280 ;
        RECT 613.830 4.000 616.210 4.280 ;
        RECT 617.050 4.000 619.890 4.280 ;
        RECT 620.730 4.000 623.570 4.280 ;
        RECT 624.410 4.000 626.790 4.280 ;
        RECT 627.630 4.000 630.470 4.280 ;
        RECT 631.310 4.000 634.150 4.280 ;
        RECT 634.990 4.000 637.370 4.280 ;
        RECT 638.210 4.000 641.050 4.280 ;
        RECT 641.890 4.000 644.730 4.280 ;
        RECT 645.570 4.000 648.410 4.280 ;
        RECT 649.250 4.000 651.630 4.280 ;
        RECT 652.470 4.000 655.310 4.280 ;
        RECT 656.150 4.000 658.990 4.280 ;
        RECT 659.830 4.000 662.210 4.280 ;
        RECT 663.050 4.000 665.890 4.280 ;
        RECT 666.730 4.000 669.570 4.280 ;
        RECT 670.410 4.000 672.790 4.280 ;
        RECT 673.630 4.000 676.470 4.280 ;
        RECT 677.310 4.000 680.150 4.280 ;
        RECT 680.990 4.000 683.370 4.280 ;
        RECT 684.210 4.000 687.050 4.280 ;
        RECT 687.890 4.000 690.730 4.280 ;
        RECT 691.570 4.000 693.950 4.280 ;
        RECT 694.790 4.000 697.630 4.280 ;
        RECT 698.470 4.000 701.310 4.280 ;
        RECT 702.150 4.000 704.990 4.280 ;
        RECT 705.830 4.000 708.210 4.280 ;
        RECT 709.050 4.000 711.890 4.280 ;
        RECT 712.730 4.000 715.570 4.280 ;
        RECT 716.410 4.000 718.790 4.280 ;
        RECT 719.630 4.000 722.470 4.280 ;
        RECT 723.310 4.000 726.150 4.280 ;
        RECT 726.990 4.000 729.370 4.280 ;
        RECT 730.210 4.000 733.050 4.280 ;
        RECT 733.890 4.000 736.730 4.280 ;
        RECT 737.570 4.000 739.950 4.280 ;
        RECT 740.790 4.000 743.630 4.280 ;
        RECT 744.470 4.000 747.310 4.280 ;
      LAYER met3 ;
        RECT 4.400 746.960 740.535 747.825 ;
        RECT 3.950 744.960 740.535 746.960 ;
        RECT 4.400 743.560 740.535 744.960 ;
        RECT 3.950 740.880 740.535 743.560 ;
        RECT 4.400 739.480 740.535 740.880 ;
        RECT 3.950 737.480 740.535 739.480 ;
        RECT 4.400 736.080 740.535 737.480 ;
        RECT 3.950 733.400 740.535 736.080 ;
        RECT 4.400 732.000 740.535 733.400 ;
        RECT 3.950 730.000 740.535 732.000 ;
        RECT 4.400 728.600 740.535 730.000 ;
        RECT 3.950 725.920 740.535 728.600 ;
        RECT 4.400 724.520 740.535 725.920 ;
        RECT 3.950 722.520 740.535 724.520 ;
        RECT 4.400 721.120 740.535 722.520 ;
        RECT 3.950 718.440 740.535 721.120 ;
        RECT 4.400 717.040 740.535 718.440 ;
        RECT 3.950 715.040 740.535 717.040 ;
        RECT 4.400 713.640 740.535 715.040 ;
        RECT 3.950 710.960 740.535 713.640 ;
        RECT 4.400 709.560 740.535 710.960 ;
        RECT 3.950 707.560 740.535 709.560 ;
        RECT 4.400 706.160 740.535 707.560 ;
        RECT 3.950 703.480 740.535 706.160 ;
        RECT 4.400 702.080 740.535 703.480 ;
        RECT 3.950 700.080 740.535 702.080 ;
        RECT 4.400 698.680 740.535 700.080 ;
        RECT 3.950 696.000 740.535 698.680 ;
        RECT 4.400 694.600 740.535 696.000 ;
        RECT 3.950 692.600 740.535 694.600 ;
        RECT 4.400 691.200 740.535 692.600 ;
        RECT 3.950 688.520 740.535 691.200 ;
        RECT 4.400 687.120 740.535 688.520 ;
        RECT 3.950 685.120 740.535 687.120 ;
        RECT 4.400 683.720 740.535 685.120 ;
        RECT 3.950 681.040 740.535 683.720 ;
        RECT 4.400 679.640 740.535 681.040 ;
        RECT 3.950 677.640 740.535 679.640 ;
        RECT 4.400 676.240 740.535 677.640 ;
        RECT 3.950 673.560 740.535 676.240 ;
        RECT 4.400 672.160 740.535 673.560 ;
        RECT 3.950 670.160 740.535 672.160 ;
        RECT 4.400 668.760 740.535 670.160 ;
        RECT 3.950 666.080 740.535 668.760 ;
        RECT 4.400 664.680 740.535 666.080 ;
        RECT 3.950 662.680 740.535 664.680 ;
        RECT 4.400 661.280 740.535 662.680 ;
        RECT 3.950 658.600 740.535 661.280 ;
        RECT 4.400 657.200 740.535 658.600 ;
        RECT 3.950 655.200 740.535 657.200 ;
        RECT 4.400 653.800 740.535 655.200 ;
        RECT 3.950 651.120 740.535 653.800 ;
        RECT 4.400 649.720 740.535 651.120 ;
        RECT 3.950 647.720 740.535 649.720 ;
        RECT 4.400 646.320 740.535 647.720 ;
        RECT 3.950 643.640 740.535 646.320 ;
        RECT 4.400 642.240 740.535 643.640 ;
        RECT 3.950 640.240 740.535 642.240 ;
        RECT 4.400 638.840 740.535 640.240 ;
        RECT 3.950 636.160 740.535 638.840 ;
        RECT 4.400 634.760 740.535 636.160 ;
        RECT 3.950 632.760 740.535 634.760 ;
        RECT 4.400 631.360 740.535 632.760 ;
        RECT 3.950 628.680 740.535 631.360 ;
        RECT 4.400 627.280 740.535 628.680 ;
        RECT 3.950 625.280 740.535 627.280 ;
        RECT 4.400 623.880 740.535 625.280 ;
        RECT 3.950 621.200 740.535 623.880 ;
        RECT 4.400 619.800 740.535 621.200 ;
        RECT 3.950 617.800 740.535 619.800 ;
        RECT 4.400 616.400 740.535 617.800 ;
        RECT 3.950 613.720 740.535 616.400 ;
        RECT 4.400 612.320 740.535 613.720 ;
        RECT 3.950 610.320 740.535 612.320 ;
        RECT 4.400 608.920 740.535 610.320 ;
        RECT 3.950 606.240 740.535 608.920 ;
        RECT 4.400 604.840 740.535 606.240 ;
        RECT 3.950 602.840 740.535 604.840 ;
        RECT 4.400 601.440 740.535 602.840 ;
        RECT 3.950 599.440 740.535 601.440 ;
        RECT 4.400 598.040 740.535 599.440 ;
        RECT 3.950 595.360 740.535 598.040 ;
        RECT 4.400 593.960 740.535 595.360 ;
        RECT 3.950 591.960 740.535 593.960 ;
        RECT 4.400 590.560 740.535 591.960 ;
        RECT 3.950 587.880 740.535 590.560 ;
        RECT 4.400 586.480 740.535 587.880 ;
        RECT 3.950 584.480 740.535 586.480 ;
        RECT 4.400 583.080 740.535 584.480 ;
        RECT 3.950 580.400 740.535 583.080 ;
        RECT 4.400 579.000 740.535 580.400 ;
        RECT 3.950 577.000 740.535 579.000 ;
        RECT 4.400 575.600 740.535 577.000 ;
        RECT 3.950 572.920 740.535 575.600 ;
        RECT 4.400 571.520 740.535 572.920 ;
        RECT 3.950 569.520 740.535 571.520 ;
        RECT 4.400 568.120 740.535 569.520 ;
        RECT 3.950 565.440 740.535 568.120 ;
        RECT 4.400 564.040 740.535 565.440 ;
        RECT 3.950 562.040 740.535 564.040 ;
        RECT 4.400 560.640 740.535 562.040 ;
        RECT 3.950 557.960 740.535 560.640 ;
        RECT 4.400 556.560 740.535 557.960 ;
        RECT 3.950 554.560 740.535 556.560 ;
        RECT 4.400 553.160 740.535 554.560 ;
        RECT 3.950 550.480 740.535 553.160 ;
        RECT 4.400 549.080 740.535 550.480 ;
        RECT 3.950 547.080 740.535 549.080 ;
        RECT 4.400 545.680 740.535 547.080 ;
        RECT 3.950 543.000 740.535 545.680 ;
        RECT 4.400 541.600 740.535 543.000 ;
        RECT 3.950 539.600 740.535 541.600 ;
        RECT 4.400 538.200 740.535 539.600 ;
        RECT 3.950 535.520 740.535 538.200 ;
        RECT 4.400 534.120 740.535 535.520 ;
        RECT 3.950 532.120 740.535 534.120 ;
        RECT 4.400 530.720 740.535 532.120 ;
        RECT 3.950 528.040 740.535 530.720 ;
        RECT 4.400 526.640 740.535 528.040 ;
        RECT 3.950 524.640 740.535 526.640 ;
        RECT 4.400 523.240 740.535 524.640 ;
        RECT 3.950 520.560 740.535 523.240 ;
        RECT 4.400 519.160 740.535 520.560 ;
        RECT 3.950 517.160 740.535 519.160 ;
        RECT 4.400 515.760 740.535 517.160 ;
        RECT 3.950 513.080 740.535 515.760 ;
        RECT 4.400 511.680 740.535 513.080 ;
        RECT 3.950 509.680 740.535 511.680 ;
        RECT 4.400 508.280 740.535 509.680 ;
        RECT 3.950 505.600 740.535 508.280 ;
        RECT 4.400 504.200 740.535 505.600 ;
        RECT 3.950 502.200 740.535 504.200 ;
        RECT 4.400 500.800 740.535 502.200 ;
        RECT 3.950 498.120 740.535 500.800 ;
        RECT 4.400 496.720 740.535 498.120 ;
        RECT 3.950 494.720 740.535 496.720 ;
        RECT 4.400 493.320 740.535 494.720 ;
        RECT 3.950 490.640 740.535 493.320 ;
        RECT 4.400 489.240 740.535 490.640 ;
        RECT 3.950 487.240 740.535 489.240 ;
        RECT 4.400 485.840 740.535 487.240 ;
        RECT 3.950 483.160 740.535 485.840 ;
        RECT 4.400 481.760 740.535 483.160 ;
        RECT 3.950 479.760 740.535 481.760 ;
        RECT 4.400 478.360 740.535 479.760 ;
        RECT 3.950 475.680 740.535 478.360 ;
        RECT 4.400 474.280 740.535 475.680 ;
        RECT 3.950 472.280 740.535 474.280 ;
        RECT 4.400 470.880 740.535 472.280 ;
        RECT 3.950 468.200 740.535 470.880 ;
        RECT 4.400 466.800 740.535 468.200 ;
        RECT 3.950 464.800 740.535 466.800 ;
        RECT 4.400 463.400 740.535 464.800 ;
        RECT 3.950 460.720 740.535 463.400 ;
        RECT 4.400 459.320 740.535 460.720 ;
        RECT 3.950 457.320 740.535 459.320 ;
        RECT 4.400 455.920 740.535 457.320 ;
        RECT 3.950 453.240 740.535 455.920 ;
        RECT 4.400 451.840 740.535 453.240 ;
        RECT 3.950 449.840 740.535 451.840 ;
        RECT 4.400 448.440 740.535 449.840 ;
        RECT 3.950 446.440 740.535 448.440 ;
        RECT 4.400 445.040 740.535 446.440 ;
        RECT 3.950 442.360 740.535 445.040 ;
        RECT 4.400 440.960 740.535 442.360 ;
        RECT 3.950 438.960 740.535 440.960 ;
        RECT 4.400 437.560 740.535 438.960 ;
        RECT 3.950 434.880 740.535 437.560 ;
        RECT 4.400 433.480 740.535 434.880 ;
        RECT 3.950 431.480 740.535 433.480 ;
        RECT 4.400 430.080 740.535 431.480 ;
        RECT 3.950 427.400 740.535 430.080 ;
        RECT 4.400 426.000 740.535 427.400 ;
        RECT 3.950 424.000 740.535 426.000 ;
        RECT 4.400 422.600 740.535 424.000 ;
        RECT 3.950 419.920 740.535 422.600 ;
        RECT 4.400 418.520 740.535 419.920 ;
        RECT 3.950 416.520 740.535 418.520 ;
        RECT 4.400 415.120 740.535 416.520 ;
        RECT 3.950 412.440 740.535 415.120 ;
        RECT 4.400 411.040 740.535 412.440 ;
        RECT 3.950 409.040 740.535 411.040 ;
        RECT 4.400 407.640 740.535 409.040 ;
        RECT 3.950 404.960 740.535 407.640 ;
        RECT 4.400 403.560 740.535 404.960 ;
        RECT 3.950 401.560 740.535 403.560 ;
        RECT 4.400 400.160 740.535 401.560 ;
        RECT 3.950 397.480 740.535 400.160 ;
        RECT 4.400 396.080 740.535 397.480 ;
        RECT 3.950 394.080 740.535 396.080 ;
        RECT 4.400 392.680 740.535 394.080 ;
        RECT 3.950 390.000 740.535 392.680 ;
        RECT 4.400 388.600 740.535 390.000 ;
        RECT 3.950 386.600 740.535 388.600 ;
        RECT 4.400 385.200 740.535 386.600 ;
        RECT 3.950 382.520 740.535 385.200 ;
        RECT 4.400 381.120 740.535 382.520 ;
        RECT 3.950 379.120 740.535 381.120 ;
        RECT 4.400 377.720 740.535 379.120 ;
        RECT 3.950 375.040 740.535 377.720 ;
        RECT 4.400 373.640 740.535 375.040 ;
        RECT 3.950 371.640 740.535 373.640 ;
        RECT 4.400 370.240 740.535 371.640 ;
        RECT 3.950 367.560 740.535 370.240 ;
        RECT 4.400 366.160 740.535 367.560 ;
        RECT 3.950 364.160 740.535 366.160 ;
        RECT 4.400 362.760 740.535 364.160 ;
        RECT 3.950 360.080 740.535 362.760 ;
        RECT 4.400 358.680 740.535 360.080 ;
        RECT 3.950 356.680 740.535 358.680 ;
        RECT 4.400 355.280 740.535 356.680 ;
        RECT 3.950 352.600 740.535 355.280 ;
        RECT 4.400 351.200 740.535 352.600 ;
        RECT 3.950 349.200 740.535 351.200 ;
        RECT 4.400 347.800 740.535 349.200 ;
        RECT 3.950 345.120 740.535 347.800 ;
        RECT 4.400 343.720 740.535 345.120 ;
        RECT 3.950 341.720 740.535 343.720 ;
        RECT 4.400 340.320 740.535 341.720 ;
        RECT 3.950 337.640 740.535 340.320 ;
        RECT 4.400 336.240 740.535 337.640 ;
        RECT 3.950 334.240 740.535 336.240 ;
        RECT 4.400 332.840 740.535 334.240 ;
        RECT 3.950 330.160 740.535 332.840 ;
        RECT 4.400 328.760 740.535 330.160 ;
        RECT 3.950 326.760 740.535 328.760 ;
        RECT 4.400 325.360 740.535 326.760 ;
        RECT 3.950 322.680 740.535 325.360 ;
        RECT 4.400 321.280 740.535 322.680 ;
        RECT 3.950 319.280 740.535 321.280 ;
        RECT 4.400 317.880 740.535 319.280 ;
        RECT 3.950 315.200 740.535 317.880 ;
        RECT 4.400 313.800 740.535 315.200 ;
        RECT 3.950 311.800 740.535 313.800 ;
        RECT 4.400 310.400 740.535 311.800 ;
        RECT 3.950 307.720 740.535 310.400 ;
        RECT 4.400 306.320 740.535 307.720 ;
        RECT 3.950 304.320 740.535 306.320 ;
        RECT 4.400 302.920 740.535 304.320 ;
        RECT 3.950 300.920 740.535 302.920 ;
        RECT 4.400 299.520 740.535 300.920 ;
        RECT 3.950 296.840 740.535 299.520 ;
        RECT 4.400 295.440 740.535 296.840 ;
        RECT 3.950 293.440 740.535 295.440 ;
        RECT 4.400 292.040 740.535 293.440 ;
        RECT 3.950 289.360 740.535 292.040 ;
        RECT 4.400 287.960 740.535 289.360 ;
        RECT 3.950 285.960 740.535 287.960 ;
        RECT 4.400 284.560 740.535 285.960 ;
        RECT 3.950 281.880 740.535 284.560 ;
        RECT 4.400 280.480 740.535 281.880 ;
        RECT 3.950 278.480 740.535 280.480 ;
        RECT 4.400 277.080 740.535 278.480 ;
        RECT 3.950 274.400 740.535 277.080 ;
        RECT 4.400 273.000 740.535 274.400 ;
        RECT 3.950 271.000 740.535 273.000 ;
        RECT 4.400 269.600 740.535 271.000 ;
        RECT 3.950 266.920 740.535 269.600 ;
        RECT 4.400 265.520 740.535 266.920 ;
        RECT 3.950 263.520 740.535 265.520 ;
        RECT 4.400 262.120 740.535 263.520 ;
        RECT 3.950 259.440 740.535 262.120 ;
        RECT 4.400 258.040 740.535 259.440 ;
        RECT 3.950 256.040 740.535 258.040 ;
        RECT 4.400 254.640 740.535 256.040 ;
        RECT 3.950 251.960 740.535 254.640 ;
        RECT 4.400 250.560 740.535 251.960 ;
        RECT 3.950 248.560 740.535 250.560 ;
        RECT 4.400 247.160 740.535 248.560 ;
        RECT 3.950 244.480 740.535 247.160 ;
        RECT 4.400 243.080 740.535 244.480 ;
        RECT 3.950 241.080 740.535 243.080 ;
        RECT 4.400 239.680 740.535 241.080 ;
        RECT 3.950 237.000 740.535 239.680 ;
        RECT 4.400 235.600 740.535 237.000 ;
        RECT 3.950 233.600 740.535 235.600 ;
        RECT 4.400 232.200 740.535 233.600 ;
        RECT 3.950 229.520 740.535 232.200 ;
        RECT 4.400 228.120 740.535 229.520 ;
        RECT 3.950 226.120 740.535 228.120 ;
        RECT 4.400 224.720 740.535 226.120 ;
        RECT 3.950 222.040 740.535 224.720 ;
        RECT 4.400 220.640 740.535 222.040 ;
        RECT 3.950 218.640 740.535 220.640 ;
        RECT 4.400 217.240 740.535 218.640 ;
        RECT 3.950 214.560 740.535 217.240 ;
        RECT 4.400 213.160 740.535 214.560 ;
        RECT 3.950 211.160 740.535 213.160 ;
        RECT 4.400 209.760 740.535 211.160 ;
        RECT 3.950 207.080 740.535 209.760 ;
        RECT 4.400 205.680 740.535 207.080 ;
        RECT 3.950 203.680 740.535 205.680 ;
        RECT 4.400 202.280 740.535 203.680 ;
        RECT 3.950 199.600 740.535 202.280 ;
        RECT 4.400 198.200 740.535 199.600 ;
        RECT 3.950 196.200 740.535 198.200 ;
        RECT 4.400 194.800 740.535 196.200 ;
        RECT 3.950 192.120 740.535 194.800 ;
        RECT 4.400 190.720 740.535 192.120 ;
        RECT 3.950 188.720 740.535 190.720 ;
        RECT 4.400 187.320 740.535 188.720 ;
        RECT 3.950 184.640 740.535 187.320 ;
        RECT 4.400 183.240 740.535 184.640 ;
        RECT 3.950 181.240 740.535 183.240 ;
        RECT 4.400 179.840 740.535 181.240 ;
        RECT 3.950 177.160 740.535 179.840 ;
        RECT 4.400 175.760 740.535 177.160 ;
        RECT 3.950 173.760 740.535 175.760 ;
        RECT 4.400 172.360 740.535 173.760 ;
        RECT 3.950 169.680 740.535 172.360 ;
        RECT 4.400 168.280 740.535 169.680 ;
        RECT 3.950 166.280 740.535 168.280 ;
        RECT 4.400 164.880 740.535 166.280 ;
        RECT 3.950 162.200 740.535 164.880 ;
        RECT 4.400 160.800 740.535 162.200 ;
        RECT 3.950 158.800 740.535 160.800 ;
        RECT 4.400 157.400 740.535 158.800 ;
        RECT 3.950 154.720 740.535 157.400 ;
        RECT 4.400 153.320 740.535 154.720 ;
        RECT 3.950 151.320 740.535 153.320 ;
        RECT 4.400 149.920 740.535 151.320 ;
        RECT 3.950 147.920 740.535 149.920 ;
        RECT 4.400 146.520 740.535 147.920 ;
        RECT 3.950 143.840 740.535 146.520 ;
        RECT 4.400 142.440 740.535 143.840 ;
        RECT 3.950 140.440 740.535 142.440 ;
        RECT 4.400 139.040 740.535 140.440 ;
        RECT 3.950 136.360 740.535 139.040 ;
        RECT 4.400 134.960 740.535 136.360 ;
        RECT 3.950 132.960 740.535 134.960 ;
        RECT 4.400 131.560 740.535 132.960 ;
        RECT 3.950 128.880 740.535 131.560 ;
        RECT 4.400 127.480 740.535 128.880 ;
        RECT 3.950 125.480 740.535 127.480 ;
        RECT 4.400 124.080 740.535 125.480 ;
        RECT 3.950 121.400 740.535 124.080 ;
        RECT 4.400 120.000 740.535 121.400 ;
        RECT 3.950 118.000 740.535 120.000 ;
        RECT 4.400 116.600 740.535 118.000 ;
        RECT 3.950 113.920 740.535 116.600 ;
        RECT 4.400 112.520 740.535 113.920 ;
        RECT 3.950 110.520 740.535 112.520 ;
        RECT 4.400 109.120 740.535 110.520 ;
        RECT 3.950 106.440 740.535 109.120 ;
        RECT 4.400 105.040 740.535 106.440 ;
        RECT 3.950 103.040 740.535 105.040 ;
        RECT 4.400 101.640 740.535 103.040 ;
        RECT 3.950 98.960 740.535 101.640 ;
        RECT 4.400 97.560 740.535 98.960 ;
        RECT 3.950 95.560 740.535 97.560 ;
        RECT 4.400 94.160 740.535 95.560 ;
        RECT 3.950 91.480 740.535 94.160 ;
        RECT 4.400 90.080 740.535 91.480 ;
        RECT 3.950 88.080 740.535 90.080 ;
        RECT 4.400 86.680 740.535 88.080 ;
        RECT 3.950 84.000 740.535 86.680 ;
        RECT 4.400 82.600 740.535 84.000 ;
        RECT 3.950 80.600 740.535 82.600 ;
        RECT 4.400 79.200 740.535 80.600 ;
        RECT 3.950 76.520 740.535 79.200 ;
        RECT 4.400 75.120 740.535 76.520 ;
        RECT 3.950 73.120 740.535 75.120 ;
        RECT 4.400 71.720 740.535 73.120 ;
        RECT 3.950 69.040 740.535 71.720 ;
        RECT 4.400 67.640 740.535 69.040 ;
        RECT 3.950 65.640 740.535 67.640 ;
        RECT 4.400 64.240 740.535 65.640 ;
        RECT 3.950 61.560 740.535 64.240 ;
        RECT 4.400 60.160 740.535 61.560 ;
        RECT 3.950 58.160 740.535 60.160 ;
        RECT 4.400 56.760 740.535 58.160 ;
        RECT 3.950 54.080 740.535 56.760 ;
        RECT 4.400 52.680 740.535 54.080 ;
        RECT 3.950 50.680 740.535 52.680 ;
        RECT 4.400 49.280 740.535 50.680 ;
        RECT 3.950 46.600 740.535 49.280 ;
        RECT 4.400 45.200 740.535 46.600 ;
        RECT 3.950 43.200 740.535 45.200 ;
        RECT 4.400 41.800 740.535 43.200 ;
        RECT 3.950 39.120 740.535 41.800 ;
        RECT 4.400 37.720 740.535 39.120 ;
        RECT 3.950 35.720 740.535 37.720 ;
        RECT 4.400 34.320 740.535 35.720 ;
        RECT 3.950 31.640 740.535 34.320 ;
        RECT 4.400 30.240 740.535 31.640 ;
        RECT 3.950 28.240 740.535 30.240 ;
        RECT 4.400 26.840 740.535 28.240 ;
        RECT 3.950 24.160 740.535 26.840 ;
        RECT 4.400 22.760 740.535 24.160 ;
        RECT 3.950 20.760 740.535 22.760 ;
        RECT 4.400 19.360 740.535 20.760 ;
        RECT 3.950 16.680 740.535 19.360 ;
        RECT 4.400 15.280 740.535 16.680 ;
        RECT 3.950 13.280 740.535 15.280 ;
        RECT 4.400 11.880 740.535 13.280 ;
        RECT 3.950 9.200 740.535 11.880 ;
        RECT 4.400 7.800 740.535 9.200 ;
        RECT 3.950 5.800 740.535 7.800 ;
        RECT 4.400 4.400 740.535 5.800 ;
        RECT 3.950 2.400 740.535 4.400 ;
        RECT 4.400 1.000 740.535 2.400 ;
        RECT 3.950 0.180 740.535 1.000 ;
      LAYER met4 ;
        RECT 3.975 737.760 732.945 738.985 ;
        RECT 3.975 10.240 20.640 737.760 ;
        RECT 23.040 737.520 97.440 737.760 ;
        RECT 23.040 10.480 23.940 737.520 ;
        RECT 26.340 10.480 27.240 737.520 ;
        RECT 29.640 10.480 30.540 737.520 ;
        RECT 32.940 10.480 97.440 737.520 ;
        RECT 23.040 10.240 97.440 10.480 ;
        RECT 99.840 737.520 174.240 737.760 ;
        RECT 99.840 10.480 100.740 737.520 ;
        RECT 103.140 10.480 104.040 737.520 ;
        RECT 106.440 10.480 107.340 737.520 ;
        RECT 109.740 10.480 174.240 737.520 ;
        RECT 99.840 10.240 174.240 10.480 ;
        RECT 176.640 737.520 251.040 737.760 ;
        RECT 176.640 10.480 177.540 737.520 ;
        RECT 179.940 10.480 180.840 737.520 ;
        RECT 183.240 10.480 184.140 737.520 ;
        RECT 186.540 10.480 251.040 737.520 ;
        RECT 176.640 10.240 251.040 10.480 ;
        RECT 253.440 737.520 327.840 737.760 ;
        RECT 253.440 10.480 254.340 737.520 ;
        RECT 256.740 10.480 257.640 737.520 ;
        RECT 260.040 10.480 260.940 737.520 ;
        RECT 263.340 10.480 327.840 737.520 ;
        RECT 253.440 10.240 327.840 10.480 ;
        RECT 330.240 737.520 404.640 737.760 ;
        RECT 330.240 10.480 331.140 737.520 ;
        RECT 333.540 10.480 334.440 737.520 ;
        RECT 336.840 10.480 337.740 737.520 ;
        RECT 340.140 10.480 404.640 737.520 ;
        RECT 330.240 10.240 404.640 10.480 ;
        RECT 407.040 737.520 481.440 737.760 ;
        RECT 407.040 10.480 407.940 737.520 ;
        RECT 410.340 10.480 411.240 737.520 ;
        RECT 413.640 10.480 414.540 737.520 ;
        RECT 416.940 10.480 481.440 737.520 ;
        RECT 407.040 10.240 481.440 10.480 ;
        RECT 483.840 737.520 558.240 737.760 ;
        RECT 483.840 10.480 484.740 737.520 ;
        RECT 487.140 10.480 488.040 737.520 ;
        RECT 490.440 10.480 491.340 737.520 ;
        RECT 493.740 10.480 558.240 737.520 ;
        RECT 483.840 10.240 558.240 10.480 ;
        RECT 560.640 737.520 635.040 737.760 ;
        RECT 560.640 10.480 561.540 737.520 ;
        RECT 563.940 10.480 564.840 737.520 ;
        RECT 567.240 10.480 568.140 737.520 ;
        RECT 570.540 10.480 635.040 737.520 ;
        RECT 560.640 10.240 635.040 10.480 ;
        RECT 637.440 737.520 711.840 737.760 ;
        RECT 637.440 10.480 638.340 737.520 ;
        RECT 640.740 10.480 641.640 737.520 ;
        RECT 644.040 10.480 644.940 737.520 ;
        RECT 647.340 10.480 711.840 737.520 ;
        RECT 637.440 10.240 711.840 10.480 ;
        RECT 714.240 737.520 732.945 737.760 ;
        RECT 714.240 10.480 715.140 737.520 ;
        RECT 717.540 10.480 718.440 737.520 ;
        RECT 720.840 10.480 721.740 737.520 ;
        RECT 724.140 10.480 732.945 737.520 ;
        RECT 714.240 10.240 732.945 10.480 ;
        RECT 3.975 0.175 732.945 10.240 ;
  END
END dcache
END LIBRARY

