VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO icache
  CLASS BLOCK ;
  FOREIGN icache ;
  ORIGIN -0.005 0.000 ;
  SIZE 678.095 BY 680.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 2.080 678.100 2.680 ;
    END
  END clk
  PIN flush_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.810 0.000 664.090 4.000 ;
    END
  END flush_in
  PIN i_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.030 0.000 0.310 4.000 ;
    END
  END i_in[0]
  PIN i_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.130 0.000 39.410 4.000 ;
    END
  END i_in[10]
  PIN i_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.810 0.000 43.090 4.000 ;
    END
  END i_in[11]
  PIN i_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.950 0.000 47.230 4.000 ;
    END
  END i_in[12]
  PIN i_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.090 0.000 51.370 4.000 ;
    END
  END i_in[13]
  PIN i_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.770 0.000 55.050 4.000 ;
    END
  END i_in[14]
  PIN i_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.910 0.000 59.190 4.000 ;
    END
  END i_in[15]
  PIN i_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.590 0.000 62.870 4.000 ;
    END
  END i_in[16]
  PIN i_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.730 0.000 67.010 4.000 ;
    END
  END i_in[17]
  PIN i_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.410 0.000 70.690 4.000 ;
    END
  END i_in[18]
  PIN i_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.550 0.000 74.830 4.000 ;
    END
  END i_in[19]
  PIN i_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.710 0.000 3.990 4.000 ;
    END
  END i_in[1]
  PIN i_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.230 0.000 78.510 4.000 ;
    END
  END i_in[20]
  PIN i_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.370 0.000 82.650 4.000 ;
    END
  END i_in[21]
  PIN i_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.050 0.000 86.330 4.000 ;
    END
  END i_in[22]
  PIN i_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.190 0.000 90.470 4.000 ;
    END
  END i_in[23]
  PIN i_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.330 0.000 94.610 4.000 ;
    END
  END i_in[24]
  PIN i_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.010 0.000 98.290 4.000 ;
    END
  END i_in[25]
  PIN i_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.150 0.000 102.430 4.000 ;
    END
  END i_in[26]
  PIN i_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.830 0.000 106.110 4.000 ;
    END
  END i_in[27]
  PIN i_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.970 0.000 110.250 4.000 ;
    END
  END i_in[28]
  PIN i_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.650 0.000 113.930 4.000 ;
    END
  END i_in[29]
  PIN i_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.850 0.000 8.130 4.000 ;
    END
  END i_in[2]
  PIN i_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.790 0.000 118.070 4.000 ;
    END
  END i_in[30]
  PIN i_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.470 0.000 121.750 4.000 ;
    END
  END i_in[31]
  PIN i_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.610 0.000 125.890 4.000 ;
    END
  END i_in[32]
  PIN i_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.290 0.000 129.570 4.000 ;
    END
  END i_in[33]
  PIN i_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.430 0.000 133.710 4.000 ;
    END
  END i_in[34]
  PIN i_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.570 0.000 137.850 4.000 ;
    END
  END i_in[35]
  PIN i_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.250 0.000 141.530 4.000 ;
    END
  END i_in[36]
  PIN i_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.390 0.000 145.670 4.000 ;
    END
  END i_in[37]
  PIN i_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.070 0.000 149.350 4.000 ;
    END
  END i_in[38]
  PIN i_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.210 0.000 153.490 4.000 ;
    END
  END i_in[39]
  PIN i_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.530 0.000 11.810 4.000 ;
    END
  END i_in[3]
  PIN i_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.890 0.000 157.170 4.000 ;
    END
  END i_in[40]
  PIN i_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.030 0.000 161.310 4.000 ;
    END
  END i_in[41]
  PIN i_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.710 0.000 164.990 4.000 ;
    END
  END i_in[42]
  PIN i_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.850 0.000 169.130 4.000 ;
    END
  END i_in[43]
  PIN i_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.530 0.000 172.810 4.000 ;
    END
  END i_in[44]
  PIN i_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.670 0.000 176.950 4.000 ;
    END
  END i_in[45]
  PIN i_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.350 0.000 180.630 4.000 ;
    END
  END i_in[46]
  PIN i_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.490 0.000 184.770 4.000 ;
    END
  END i_in[47]
  PIN i_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.630 0.000 188.910 4.000 ;
    END
  END i_in[48]
  PIN i_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.310 0.000 192.590 4.000 ;
    END
  END i_in[49]
  PIN i_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.670 0.000 15.950 4.000 ;
    END
  END i_in[4]
  PIN i_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.450 0.000 196.730 4.000 ;
    END
  END i_in[50]
  PIN i_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.130 0.000 200.410 4.000 ;
    END
  END i_in[51]
  PIN i_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.270 0.000 204.550 4.000 ;
    END
  END i_in[52]
  PIN i_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.950 0.000 208.230 4.000 ;
    END
  END i_in[53]
  PIN i_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.090 0.000 212.370 4.000 ;
    END
  END i_in[54]
  PIN i_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.770 0.000 216.050 4.000 ;
    END
  END i_in[55]
  PIN i_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.910 0.000 220.190 4.000 ;
    END
  END i_in[56]
  PIN i_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.590 0.000 223.870 4.000 ;
    END
  END i_in[57]
  PIN i_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.730 0.000 228.010 4.000 ;
    END
  END i_in[58]
  PIN i_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.870 0.000 232.150 4.000 ;
    END
  END i_in[59]
  PIN i_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.350 0.000 19.630 4.000 ;
    END
  END i_in[5]
  PIN i_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.550 0.000 235.830 4.000 ;
    END
  END i_in[60]
  PIN i_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.690 0.000 239.970 4.000 ;
    END
  END i_in[61]
  PIN i_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.370 0.000 243.650 4.000 ;
    END
  END i_in[62]
  PIN i_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.510 0.000 247.790 4.000 ;
    END
  END i_in[63]
  PIN i_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.190 0.000 251.470 4.000 ;
    END
  END i_in[64]
  PIN i_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.330 0.000 255.610 4.000 ;
    END
  END i_in[65]
  PIN i_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.010 0.000 259.290 4.000 ;
    END
  END i_in[66]
  PIN i_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.150 0.000 263.430 4.000 ;
    END
  END i_in[67]
  PIN i_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.830 0.000 267.110 4.000 ;
    END
  END i_in[68]
  PIN i_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.970 0.000 271.250 4.000 ;
    END
  END i_in[69]
  PIN i_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.490 0.000 23.770 4.000 ;
    END
  END i_in[6]
  PIN i_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.170 0.000 27.450 4.000 ;
    END
  END i_in[7]
  PIN i_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.310 0.000 31.590 4.000 ;
    END
  END i_in[8]
  PIN i_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.990 0.000 35.270 4.000 ;
    END
  END i_in[9]
  PIN i_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.110 0.000 275.390 4.000 ;
    END
  END i_out[0]
  PIN i_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.210 0.000 314.490 4.000 ;
    END
  END i_out[10]
  PIN i_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.350 0.000 318.630 4.000 ;
    END
  END i_out[11]
  PIN i_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.030 0.000 322.310 4.000 ;
    END
  END i_out[12]
  PIN i_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.170 0.000 326.450 4.000 ;
    END
  END i_out[13]
  PIN i_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.850 0.000 330.130 4.000 ;
    END
  END i_out[14]
  PIN i_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.990 0.000 334.270 4.000 ;
    END
  END i_out[15]
  PIN i_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.670 0.000 337.950 4.000 ;
    END
  END i_out[16]
  PIN i_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.810 0.000 342.090 4.000 ;
    END
  END i_out[17]
  PIN i_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.490 0.000 345.770 4.000 ;
    END
  END i_out[18]
  PIN i_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.630 0.000 349.910 4.000 ;
    END
  END i_out[19]
  PIN i_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.790 0.000 279.070 4.000 ;
    END
  END i_out[1]
  PIN i_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.310 0.000 353.590 4.000 ;
    END
  END i_out[20]
  PIN i_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.450 0.000 357.730 4.000 ;
    END
  END i_out[21]
  PIN i_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.130 0.000 361.410 4.000 ;
    END
  END i_out[22]
  PIN i_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.270 0.000 365.550 4.000 ;
    END
  END i_out[23]
  PIN i_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.410 0.000 369.690 4.000 ;
    END
  END i_out[24]
  PIN i_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.090 0.000 373.370 4.000 ;
    END
  END i_out[25]
  PIN i_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.230 0.000 377.510 4.000 ;
    END
  END i_out[26]
  PIN i_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.910 0.000 381.190 4.000 ;
    END
  END i_out[27]
  PIN i_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.050 0.000 385.330 4.000 ;
    END
  END i_out[28]
  PIN i_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.730 0.000 389.010 4.000 ;
    END
  END i_out[29]
  PIN i_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.930 0.000 283.210 4.000 ;
    END
  END i_out[2]
  PIN i_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.870 0.000 393.150 4.000 ;
    END
  END i_out[30]
  PIN i_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.550 0.000 396.830 4.000 ;
    END
  END i_out[31]
  PIN i_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.690 0.000 400.970 4.000 ;
    END
  END i_out[32]
  PIN i_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.370 0.000 404.650 4.000 ;
    END
  END i_out[33]
  PIN i_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.510 0.000 408.790 4.000 ;
    END
  END i_out[34]
  PIN i_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.650 0.000 412.930 4.000 ;
    END
  END i_out[35]
  PIN i_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.330 0.000 416.610 4.000 ;
    END
  END i_out[36]
  PIN i_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.470 0.000 420.750 4.000 ;
    END
  END i_out[37]
  PIN i_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.150 0.000 424.430 4.000 ;
    END
  END i_out[38]
  PIN i_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.290 0.000 428.570 4.000 ;
    END
  END i_out[39]
  PIN i_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.610 0.000 286.890 4.000 ;
    END
  END i_out[3]
  PIN i_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.970 0.000 432.250 4.000 ;
    END
  END i_out[40]
  PIN i_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.110 0.000 436.390 4.000 ;
    END
  END i_out[41]
  PIN i_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.790 0.000 440.070 4.000 ;
    END
  END i_out[42]
  PIN i_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.930 0.000 444.210 4.000 ;
    END
  END i_out[43]
  PIN i_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.610 0.000 447.890 4.000 ;
    END
  END i_out[44]
  PIN i_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.750 0.000 452.030 4.000 ;
    END
  END i_out[45]
  PIN i_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.890 0.000 456.170 4.000 ;
    END
  END i_out[46]
  PIN i_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.570 0.000 459.850 4.000 ;
    END
  END i_out[47]
  PIN i_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.710 0.000 463.990 4.000 ;
    END
  END i_out[48]
  PIN i_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.390 0.000 467.670 4.000 ;
    END
  END i_out[49]
  PIN i_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.750 0.000 291.030 4.000 ;
    END
  END i_out[4]
  PIN i_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.530 0.000 471.810 4.000 ;
    END
  END i_out[50]
  PIN i_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.210 0.000 475.490 4.000 ;
    END
  END i_out[51]
  PIN i_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.350 0.000 479.630 4.000 ;
    END
  END i_out[52]
  PIN i_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.030 0.000 483.310 4.000 ;
    END
  END i_out[53]
  PIN i_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.170 0.000 487.450 4.000 ;
    END
  END i_out[54]
  PIN i_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.850 0.000 491.130 4.000 ;
    END
  END i_out[55]
  PIN i_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.990 0.000 495.270 4.000 ;
    END
  END i_out[56]
  PIN i_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.130 0.000 499.410 4.000 ;
    END
  END i_out[57]
  PIN i_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.810 0.000 503.090 4.000 ;
    END
  END i_out[58]
  PIN i_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.950 0.000 507.230 4.000 ;
    END
  END i_out[59]
  PIN i_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.430 0.000 294.710 4.000 ;
    END
  END i_out[5]
  PIN i_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.630 0.000 510.910 4.000 ;
    END
  END i_out[60]
  PIN i_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.770 0.000 515.050 4.000 ;
    END
  END i_out[61]
  PIN i_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.450 0.000 518.730 4.000 ;
    END
  END i_out[62]
  PIN i_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.590 0.000 522.870 4.000 ;
    END
  END i_out[63]
  PIN i_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.270 0.000 526.550 4.000 ;
    END
  END i_out[64]
  PIN i_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.410 0.000 530.690 4.000 ;
    END
  END i_out[65]
  PIN i_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.090 0.000 534.370 4.000 ;
    END
  END i_out[66]
  PIN i_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.230 0.000 538.510 4.000 ;
    END
  END i_out[67]
  PIN i_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.910 0.000 542.190 4.000 ;
    END
  END i_out[68]
  PIN i_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.050 0.000 546.330 4.000 ;
    END
  END i_out[69]
  PIN i_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.570 0.000 298.850 4.000 ;
    END
  END i_out[6]
  PIN i_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.190 0.000 550.470 4.000 ;
    END
  END i_out[70]
  PIN i_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.870 0.000 554.150 4.000 ;
    END
  END i_out[71]
  PIN i_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.010 0.000 558.290 4.000 ;
    END
  END i_out[72]
  PIN i_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.690 0.000 561.970 4.000 ;
    END
  END i_out[73]
  PIN i_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.830 0.000 566.110 4.000 ;
    END
  END i_out[74]
  PIN i_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.510 0.000 569.790 4.000 ;
    END
  END i_out[75]
  PIN i_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.650 0.000 573.930 4.000 ;
    END
  END i_out[76]
  PIN i_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.330 0.000 577.610 4.000 ;
    END
  END i_out[77]
  PIN i_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.470 0.000 581.750 4.000 ;
    END
  END i_out[78]
  PIN i_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.150 0.000 585.430 4.000 ;
    END
  END i_out[79]
  PIN i_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.250 0.000 302.530 4.000 ;
    END
  END i_out[7]
  PIN i_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.290 0.000 589.570 4.000 ;
    END
  END i_out[80]
  PIN i_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.430 0.000 593.710 4.000 ;
    END
  END i_out[81]
  PIN i_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.110 0.000 597.390 4.000 ;
    END
  END i_out[82]
  PIN i_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.250 0.000 601.530 4.000 ;
    END
  END i_out[83]
  PIN i_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.930 0.000 605.210 4.000 ;
    END
  END i_out[84]
  PIN i_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.070 0.000 609.350 4.000 ;
    END
  END i_out[85]
  PIN i_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.750 0.000 613.030 4.000 ;
    END
  END i_out[86]
  PIN i_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.890 0.000 617.170 4.000 ;
    END
  END i_out[87]
  PIN i_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.570 0.000 620.850 4.000 ;
    END
  END i_out[88]
  PIN i_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.710 0.000 624.990 4.000 ;
    END
  END i_out[89]
  PIN i_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.390 0.000 306.670 4.000 ;
    END
  END i_out[8]
  PIN i_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.390 0.000 628.670 4.000 ;
    END
  END i_out[90]
  PIN i_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.530 0.000 632.810 4.000 ;
    END
  END i_out[91]
  PIN i_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.670 0.000 636.950 4.000 ;
    END
  END i_out[92]
  PIN i_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.350 0.000 640.630 4.000 ;
    END
  END i_out[93]
  PIN i_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.490 0.000 644.770 4.000 ;
    END
  END i_out[94]
  PIN i_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.170 0.000 648.450 4.000 ;
    END
  END i_out[95]
  PIN i_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.310 0.000 652.590 4.000 ;
    END
  END i_out[96]
  PIN i_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.990 0.000 656.270 4.000 ;
    END
  END i_out[97]
  PIN i_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.130 0.000 660.410 4.000 ;
    END
  END i_out[98]
  PIN i_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.070 0.000 310.350 4.000 ;
    END
  END i_out[9]
  PIN inval_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.950 0.000 668.230 4.000 ;
    END
  END inval_in
  PIN m_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 12.280 678.100 12.880 ;
    END
  END m_in[0]
  PIN m_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 522.960 678.100 523.560 ;
    END
  END m_in[100]
  PIN m_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 528.400 678.100 529.000 ;
    END
  END m_in[101]
  PIN m_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 533.160 678.100 533.760 ;
    END
  END m_in[102]
  PIN m_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 538.600 678.100 539.200 ;
    END
  END m_in[103]
  PIN m_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 543.360 678.100 543.960 ;
    END
  END m_in[104]
  PIN m_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 548.800 678.100 549.400 ;
    END
  END m_in[105]
  PIN m_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 554.240 678.100 554.840 ;
    END
  END m_in[106]
  PIN m_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 559.000 678.100 559.600 ;
    END
  END m_in[107]
  PIN m_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 564.440 678.100 565.040 ;
    END
  END m_in[108]
  PIN m_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 569.200 678.100 569.800 ;
    END
  END m_in[109]
  PIN m_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 63.280 678.100 63.880 ;
    END
  END m_in[10]
  PIN m_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 574.640 678.100 575.240 ;
    END
  END m_in[110]
  PIN m_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 579.400 678.100 580.000 ;
    END
  END m_in[111]
  PIN m_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 584.840 678.100 585.440 ;
    END
  END m_in[112]
  PIN m_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 589.600 678.100 590.200 ;
    END
  END m_in[113]
  PIN m_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 595.040 678.100 595.640 ;
    END
  END m_in[114]
  PIN m_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 599.800 678.100 600.400 ;
    END
  END m_in[115]
  PIN m_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 605.240 678.100 605.840 ;
    END
  END m_in[116]
  PIN m_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 610.000 678.100 610.600 ;
    END
  END m_in[117]
  PIN m_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 615.440 678.100 616.040 ;
    END
  END m_in[118]
  PIN m_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 620.200 678.100 620.800 ;
    END
  END m_in[119]
  PIN m_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 68.040 678.100 68.640 ;
    END
  END m_in[11]
  PIN m_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 625.640 678.100 626.240 ;
    END
  END m_in[120]
  PIN m_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 630.400 678.100 631.000 ;
    END
  END m_in[121]
  PIN m_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 635.840 678.100 636.440 ;
    END
  END m_in[122]
  PIN m_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 640.600 678.100 641.200 ;
    END
  END m_in[123]
  PIN m_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 646.040 678.100 646.640 ;
    END
  END m_in[124]
  PIN m_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 650.800 678.100 651.400 ;
    END
  END m_in[125]
  PIN m_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 656.240 678.100 656.840 ;
    END
  END m_in[126]
  PIN m_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 661.000 678.100 661.600 ;
    END
  END m_in[127]
  PIN m_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 666.440 678.100 667.040 ;
    END
  END m_in[128]
  PIN m_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 671.200 678.100 671.800 ;
    END
  END m_in[129]
  PIN m_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 73.480 678.100 74.080 ;
    END
  END m_in[12]
  PIN m_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 676.640 678.100 677.240 ;
    END
  END m_in[130]
  PIN m_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 78.240 678.100 78.840 ;
    END
  END m_in[13]
  PIN m_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 83.680 678.100 84.280 ;
    END
  END m_in[14]
  PIN m_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 88.440 678.100 89.040 ;
    END
  END m_in[15]
  PIN m_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 93.880 678.100 94.480 ;
    END
  END m_in[16]
  PIN m_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 98.640 678.100 99.240 ;
    END
  END m_in[17]
  PIN m_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 104.080 678.100 104.680 ;
    END
  END m_in[18]
  PIN m_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 108.840 678.100 109.440 ;
    END
  END m_in[19]
  PIN m_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 17.040 678.100 17.640 ;
    END
  END m_in[1]
  PIN m_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 114.280 678.100 114.880 ;
    END
  END m_in[20]
  PIN m_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 119.040 678.100 119.640 ;
    END
  END m_in[21]
  PIN m_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 124.480 678.100 125.080 ;
    END
  END m_in[22]
  PIN m_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 129.240 678.100 129.840 ;
    END
  END m_in[23]
  PIN m_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 134.680 678.100 135.280 ;
    END
  END m_in[24]
  PIN m_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 140.120 678.100 140.720 ;
    END
  END m_in[25]
  PIN m_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 144.880 678.100 145.480 ;
    END
  END m_in[26]
  PIN m_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 150.320 678.100 150.920 ;
    END
  END m_in[27]
  PIN m_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 155.080 678.100 155.680 ;
    END
  END m_in[28]
  PIN m_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 160.520 678.100 161.120 ;
    END
  END m_in[29]
  PIN m_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 22.480 678.100 23.080 ;
    END
  END m_in[2]
  PIN m_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 165.280 678.100 165.880 ;
    END
  END m_in[30]
  PIN m_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 170.720 678.100 171.320 ;
    END
  END m_in[31]
  PIN m_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 175.480 678.100 176.080 ;
    END
  END m_in[32]
  PIN m_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 180.920 678.100 181.520 ;
    END
  END m_in[33]
  PIN m_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 185.680 678.100 186.280 ;
    END
  END m_in[34]
  PIN m_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 191.120 678.100 191.720 ;
    END
  END m_in[35]
  PIN m_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 195.880 678.100 196.480 ;
    END
  END m_in[36]
  PIN m_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 201.320 678.100 201.920 ;
    END
  END m_in[37]
  PIN m_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 206.080 678.100 206.680 ;
    END
  END m_in[38]
  PIN m_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 211.520 678.100 212.120 ;
    END
  END m_in[39]
  PIN m_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 27.240 678.100 27.840 ;
    END
  END m_in[3]
  PIN m_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 216.280 678.100 216.880 ;
    END
  END m_in[40]
  PIN m_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 221.720 678.100 222.320 ;
    END
  END m_in[41]
  PIN m_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 226.480 678.100 227.080 ;
    END
  END m_in[42]
  PIN m_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 231.920 678.100 232.520 ;
    END
  END m_in[43]
  PIN m_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 236.680 678.100 237.280 ;
    END
  END m_in[44]
  PIN m_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 242.120 678.100 242.720 ;
    END
  END m_in[45]
  PIN m_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 246.880 678.100 247.480 ;
    END
  END m_in[46]
  PIN m_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 252.320 678.100 252.920 ;
    END
  END m_in[47]
  PIN m_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 257.080 678.100 257.680 ;
    END
  END m_in[48]
  PIN m_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 262.520 678.100 263.120 ;
    END
  END m_in[49]
  PIN m_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 32.680 678.100 33.280 ;
    END
  END m_in[4]
  PIN m_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 267.280 678.100 267.880 ;
    END
  END m_in[50]
  PIN m_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 272.720 678.100 273.320 ;
    END
  END m_in[51]
  PIN m_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 278.160 678.100 278.760 ;
    END
  END m_in[52]
  PIN m_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 282.920 678.100 283.520 ;
    END
  END m_in[53]
  PIN m_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 288.360 678.100 288.960 ;
    END
  END m_in[54]
  PIN m_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 293.120 678.100 293.720 ;
    END
  END m_in[55]
  PIN m_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 298.560 678.100 299.160 ;
    END
  END m_in[56]
  PIN m_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 303.320 678.100 303.920 ;
    END
  END m_in[57]
  PIN m_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 308.760 678.100 309.360 ;
    END
  END m_in[58]
  PIN m_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 313.520 678.100 314.120 ;
    END
  END m_in[59]
  PIN m_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 37.440 678.100 38.040 ;
    END
  END m_in[5]
  PIN m_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 318.960 678.100 319.560 ;
    END
  END m_in[60]
  PIN m_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 323.720 678.100 324.320 ;
    END
  END m_in[61]
  PIN m_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 329.160 678.100 329.760 ;
    END
  END m_in[62]
  PIN m_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 333.920 678.100 334.520 ;
    END
  END m_in[63]
  PIN m_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 339.360 678.100 339.960 ;
    END
  END m_in[64]
  PIN m_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 344.120 678.100 344.720 ;
    END
  END m_in[65]
  PIN m_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 349.560 678.100 350.160 ;
    END
  END m_in[66]
  PIN m_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 354.320 678.100 354.920 ;
    END
  END m_in[67]
  PIN m_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 359.760 678.100 360.360 ;
    END
  END m_in[68]
  PIN m_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 364.520 678.100 365.120 ;
    END
  END m_in[69]
  PIN m_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 42.880 678.100 43.480 ;
    END
  END m_in[6]
  PIN m_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 369.960 678.100 370.560 ;
    END
  END m_in[70]
  PIN m_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 374.720 678.100 375.320 ;
    END
  END m_in[71]
  PIN m_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 380.160 678.100 380.760 ;
    END
  END m_in[72]
  PIN m_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 384.920 678.100 385.520 ;
    END
  END m_in[73]
  PIN m_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 390.360 678.100 390.960 ;
    END
  END m_in[74]
  PIN m_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 395.120 678.100 395.720 ;
    END
  END m_in[75]
  PIN m_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 400.560 678.100 401.160 ;
    END
  END m_in[76]
  PIN m_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 405.320 678.100 405.920 ;
    END
  END m_in[77]
  PIN m_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 410.760 678.100 411.360 ;
    END
  END m_in[78]
  PIN m_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 416.200 678.100 416.800 ;
    END
  END m_in[79]
  PIN m_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 47.640 678.100 48.240 ;
    END
  END m_in[7]
  PIN m_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 420.960 678.100 421.560 ;
    END
  END m_in[80]
  PIN m_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 426.400 678.100 427.000 ;
    END
  END m_in[81]
  PIN m_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 431.160 678.100 431.760 ;
    END
  END m_in[82]
  PIN m_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 436.600 678.100 437.200 ;
    END
  END m_in[83]
  PIN m_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 441.360 678.100 441.960 ;
    END
  END m_in[84]
  PIN m_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 446.800 678.100 447.400 ;
    END
  END m_in[85]
  PIN m_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 451.560 678.100 452.160 ;
    END
  END m_in[86]
  PIN m_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 457.000 678.100 457.600 ;
    END
  END m_in[87]
  PIN m_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 461.760 678.100 462.360 ;
    END
  END m_in[88]
  PIN m_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 467.200 678.100 467.800 ;
    END
  END m_in[89]
  PIN m_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 53.080 678.100 53.680 ;
    END
  END m_in[8]
  PIN m_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 471.960 678.100 472.560 ;
    END
  END m_in[90]
  PIN m_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 477.400 678.100 478.000 ;
    END
  END m_in[91]
  PIN m_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 482.160 678.100 482.760 ;
    END
  END m_in[92]
  PIN m_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 487.600 678.100 488.200 ;
    END
  END m_in[93]
  PIN m_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 492.360 678.100 492.960 ;
    END
  END m_in[94]
  PIN m_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 497.800 678.100 498.400 ;
    END
  END m_in[95]
  PIN m_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 502.560 678.100 503.160 ;
    END
  END m_in[96]
  PIN m_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 508.000 678.100 508.600 ;
    END
  END m_in[97]
  PIN m_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 512.760 678.100 513.360 ;
    END
  END m_in[98]
  PIN m_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 518.200 678.100 518.800 ;
    END
  END m_in[99]
  PIN m_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 57.840 678.100 58.440 ;
    END
  END m_in[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 674.100 6.840 678.100 7.440 ;
    END
  END rst
  PIN stall_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.630 0.000 671.910 4.000 ;
    END
  END stall_in
  PIN stall_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.770 0.000 676.050 4.000 ;
    END
  END stall_out
  PIN wishbone_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.030 676.000 0.310 680.000 ;
    END
  END wishbone_in[0]
  PIN wishbone_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.130 676.000 39.410 680.000 ;
    END
  END wishbone_in[10]
  PIN wishbone_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.810 676.000 43.090 680.000 ;
    END
  END wishbone_in[11]
  PIN wishbone_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.950 676.000 47.230 680.000 ;
    END
  END wishbone_in[12]
  PIN wishbone_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.090 676.000 51.370 680.000 ;
    END
  END wishbone_in[13]
  PIN wishbone_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.770 676.000 55.050 680.000 ;
    END
  END wishbone_in[14]
  PIN wishbone_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.910 676.000 59.190 680.000 ;
    END
  END wishbone_in[15]
  PIN wishbone_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.590 676.000 62.870 680.000 ;
    END
  END wishbone_in[16]
  PIN wishbone_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.730 676.000 67.010 680.000 ;
    END
  END wishbone_in[17]
  PIN wishbone_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.410 676.000 70.690 680.000 ;
    END
  END wishbone_in[18]
  PIN wishbone_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.550 676.000 74.830 680.000 ;
    END
  END wishbone_in[19]
  PIN wishbone_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.710 676.000 3.990 680.000 ;
    END
  END wishbone_in[1]
  PIN wishbone_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.230 676.000 78.510 680.000 ;
    END
  END wishbone_in[20]
  PIN wishbone_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.370 676.000 82.650 680.000 ;
    END
  END wishbone_in[21]
  PIN wishbone_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.050 676.000 86.330 680.000 ;
    END
  END wishbone_in[22]
  PIN wishbone_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.190 676.000 90.470 680.000 ;
    END
  END wishbone_in[23]
  PIN wishbone_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.330 676.000 94.610 680.000 ;
    END
  END wishbone_in[24]
  PIN wishbone_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.010 676.000 98.290 680.000 ;
    END
  END wishbone_in[25]
  PIN wishbone_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.150 676.000 102.430 680.000 ;
    END
  END wishbone_in[26]
  PIN wishbone_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.830 676.000 106.110 680.000 ;
    END
  END wishbone_in[27]
  PIN wishbone_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.970 676.000 110.250 680.000 ;
    END
  END wishbone_in[28]
  PIN wishbone_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.650 676.000 113.930 680.000 ;
    END
  END wishbone_in[29]
  PIN wishbone_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.850 676.000 8.130 680.000 ;
    END
  END wishbone_in[2]
  PIN wishbone_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.790 676.000 118.070 680.000 ;
    END
  END wishbone_in[30]
  PIN wishbone_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.470 676.000 121.750 680.000 ;
    END
  END wishbone_in[31]
  PIN wishbone_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.610 676.000 125.890 680.000 ;
    END
  END wishbone_in[32]
  PIN wishbone_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.290 676.000 129.570 680.000 ;
    END
  END wishbone_in[33]
  PIN wishbone_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.430 676.000 133.710 680.000 ;
    END
  END wishbone_in[34]
  PIN wishbone_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.570 676.000 137.850 680.000 ;
    END
  END wishbone_in[35]
  PIN wishbone_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.250 676.000 141.530 680.000 ;
    END
  END wishbone_in[36]
  PIN wishbone_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.390 676.000 145.670 680.000 ;
    END
  END wishbone_in[37]
  PIN wishbone_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.070 676.000 149.350 680.000 ;
    END
  END wishbone_in[38]
  PIN wishbone_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.210 676.000 153.490 680.000 ;
    END
  END wishbone_in[39]
  PIN wishbone_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.530 676.000 11.810 680.000 ;
    END
  END wishbone_in[3]
  PIN wishbone_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.890 676.000 157.170 680.000 ;
    END
  END wishbone_in[40]
  PIN wishbone_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.030 676.000 161.310 680.000 ;
    END
  END wishbone_in[41]
  PIN wishbone_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.710 676.000 164.990 680.000 ;
    END
  END wishbone_in[42]
  PIN wishbone_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.850 676.000 169.130 680.000 ;
    END
  END wishbone_in[43]
  PIN wishbone_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.530 676.000 172.810 680.000 ;
    END
  END wishbone_in[44]
  PIN wishbone_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.670 676.000 176.950 680.000 ;
    END
  END wishbone_in[45]
  PIN wishbone_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.350 676.000 180.630 680.000 ;
    END
  END wishbone_in[46]
  PIN wishbone_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.490 676.000 184.770 680.000 ;
    END
  END wishbone_in[47]
  PIN wishbone_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.630 676.000 188.910 680.000 ;
    END
  END wishbone_in[48]
  PIN wishbone_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.310 676.000 192.590 680.000 ;
    END
  END wishbone_in[49]
  PIN wishbone_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.670 676.000 15.950 680.000 ;
    END
  END wishbone_in[4]
  PIN wishbone_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.450 676.000 196.730 680.000 ;
    END
  END wishbone_in[50]
  PIN wishbone_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.130 676.000 200.410 680.000 ;
    END
  END wishbone_in[51]
  PIN wishbone_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.270 676.000 204.550 680.000 ;
    END
  END wishbone_in[52]
  PIN wishbone_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.950 676.000 208.230 680.000 ;
    END
  END wishbone_in[53]
  PIN wishbone_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.090 676.000 212.370 680.000 ;
    END
  END wishbone_in[54]
  PIN wishbone_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.770 676.000 216.050 680.000 ;
    END
  END wishbone_in[55]
  PIN wishbone_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.910 676.000 220.190 680.000 ;
    END
  END wishbone_in[56]
  PIN wishbone_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.590 676.000 223.870 680.000 ;
    END
  END wishbone_in[57]
  PIN wishbone_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.730 676.000 228.010 680.000 ;
    END
  END wishbone_in[58]
  PIN wishbone_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.870 676.000 232.150 680.000 ;
    END
  END wishbone_in[59]
  PIN wishbone_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.350 676.000 19.630 680.000 ;
    END
  END wishbone_in[5]
  PIN wishbone_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.550 676.000 235.830 680.000 ;
    END
  END wishbone_in[60]
  PIN wishbone_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.690 676.000 239.970 680.000 ;
    END
  END wishbone_in[61]
  PIN wishbone_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.370 676.000 243.650 680.000 ;
    END
  END wishbone_in[62]
  PIN wishbone_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.510 676.000 247.790 680.000 ;
    END
  END wishbone_in[63]
  PIN wishbone_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.190 676.000 251.470 680.000 ;
    END
  END wishbone_in[64]
  PIN wishbone_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.330 676.000 255.610 680.000 ;
    END
  END wishbone_in[65]
  PIN wishbone_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.490 676.000 23.770 680.000 ;
    END
  END wishbone_in[6]
  PIN wishbone_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.170 676.000 27.450 680.000 ;
    END
  END wishbone_in[7]
  PIN wishbone_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.310 676.000 31.590 680.000 ;
    END
  END wishbone_in[8]
  PIN wishbone_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.990 676.000 35.270 680.000 ;
    END
  END wishbone_in[9]
  PIN wishbone_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.010 676.000 259.290 680.000 ;
    END
  END wishbone_out[0]
  PIN wishbone_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.310 676.000 652.590 680.000 ;
    END
  END wishbone_out[100]
  PIN wishbone_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.990 676.000 656.270 680.000 ;
    END
  END wishbone_out[101]
  PIN wishbone_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.130 676.000 660.410 680.000 ;
    END
  END wishbone_out[102]
  PIN wishbone_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.810 676.000 664.090 680.000 ;
    END
  END wishbone_out[103]
  PIN wishbone_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.950 676.000 668.230 680.000 ;
    END
  END wishbone_out[104]
  PIN wishbone_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.630 676.000 671.910 680.000 ;
    END
  END wishbone_out[105]
  PIN wishbone_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.770 676.000 676.050 680.000 ;
    END
  END wishbone_out[106]
  PIN wishbone_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.570 676.000 298.850 680.000 ;
    END
  END wishbone_out[10]
  PIN wishbone_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.250 676.000 302.530 680.000 ;
    END
  END wishbone_out[11]
  PIN wishbone_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.390 676.000 306.670 680.000 ;
    END
  END wishbone_out[12]
  PIN wishbone_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.070 676.000 310.350 680.000 ;
    END
  END wishbone_out[13]
  PIN wishbone_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.210 676.000 314.490 680.000 ;
    END
  END wishbone_out[14]
  PIN wishbone_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.350 676.000 318.630 680.000 ;
    END
  END wishbone_out[15]
  PIN wishbone_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.030 676.000 322.310 680.000 ;
    END
  END wishbone_out[16]
  PIN wishbone_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.170 676.000 326.450 680.000 ;
    END
  END wishbone_out[17]
  PIN wishbone_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.850 676.000 330.130 680.000 ;
    END
  END wishbone_out[18]
  PIN wishbone_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.990 676.000 334.270 680.000 ;
    END
  END wishbone_out[19]
  PIN wishbone_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.150 676.000 263.430 680.000 ;
    END
  END wishbone_out[1]
  PIN wishbone_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.670 676.000 337.950 680.000 ;
    END
  END wishbone_out[20]
  PIN wishbone_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.810 676.000 342.090 680.000 ;
    END
  END wishbone_out[21]
  PIN wishbone_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.490 676.000 345.770 680.000 ;
    END
  END wishbone_out[22]
  PIN wishbone_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.630 676.000 349.910 680.000 ;
    END
  END wishbone_out[23]
  PIN wishbone_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.310 676.000 353.590 680.000 ;
    END
  END wishbone_out[24]
  PIN wishbone_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.450 676.000 357.730 680.000 ;
    END
  END wishbone_out[25]
  PIN wishbone_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.130 676.000 361.410 680.000 ;
    END
  END wishbone_out[26]
  PIN wishbone_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.270 676.000 365.550 680.000 ;
    END
  END wishbone_out[27]
  PIN wishbone_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.410 676.000 369.690 680.000 ;
    END
  END wishbone_out[28]
  PIN wishbone_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.090 676.000 373.370 680.000 ;
    END
  END wishbone_out[29]
  PIN wishbone_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.830 676.000 267.110 680.000 ;
    END
  END wishbone_out[2]
  PIN wishbone_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.230 676.000 377.510 680.000 ;
    END
  END wishbone_out[30]
  PIN wishbone_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.910 676.000 381.190 680.000 ;
    END
  END wishbone_out[31]
  PIN wishbone_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.050 676.000 385.330 680.000 ;
    END
  END wishbone_out[32]
  PIN wishbone_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.730 676.000 389.010 680.000 ;
    END
  END wishbone_out[33]
  PIN wishbone_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.870 676.000 393.150 680.000 ;
    END
  END wishbone_out[34]
  PIN wishbone_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.550 676.000 396.830 680.000 ;
    END
  END wishbone_out[35]
  PIN wishbone_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.690 676.000 400.970 680.000 ;
    END
  END wishbone_out[36]
  PIN wishbone_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.370 676.000 404.650 680.000 ;
    END
  END wishbone_out[37]
  PIN wishbone_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.510 676.000 408.790 680.000 ;
    END
  END wishbone_out[38]
  PIN wishbone_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.650 676.000 412.930 680.000 ;
    END
  END wishbone_out[39]
  PIN wishbone_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.970 676.000 271.250 680.000 ;
    END
  END wishbone_out[3]
  PIN wishbone_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.330 676.000 416.610 680.000 ;
    END
  END wishbone_out[40]
  PIN wishbone_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.470 676.000 420.750 680.000 ;
    END
  END wishbone_out[41]
  PIN wishbone_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.150 676.000 424.430 680.000 ;
    END
  END wishbone_out[42]
  PIN wishbone_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.290 676.000 428.570 680.000 ;
    END
  END wishbone_out[43]
  PIN wishbone_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.970 676.000 432.250 680.000 ;
    END
  END wishbone_out[44]
  PIN wishbone_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.110 676.000 436.390 680.000 ;
    END
  END wishbone_out[45]
  PIN wishbone_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.790 676.000 440.070 680.000 ;
    END
  END wishbone_out[46]
  PIN wishbone_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.930 676.000 444.210 680.000 ;
    END
  END wishbone_out[47]
  PIN wishbone_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.610 676.000 447.890 680.000 ;
    END
  END wishbone_out[48]
  PIN wishbone_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.750 676.000 452.030 680.000 ;
    END
  END wishbone_out[49]
  PIN wishbone_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.110 676.000 275.390 680.000 ;
    END
  END wishbone_out[4]
  PIN wishbone_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.890 676.000 456.170 680.000 ;
    END
  END wishbone_out[50]
  PIN wishbone_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.570 676.000 459.850 680.000 ;
    END
  END wishbone_out[51]
  PIN wishbone_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.710 676.000 463.990 680.000 ;
    END
  END wishbone_out[52]
  PIN wishbone_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.390 676.000 467.670 680.000 ;
    END
  END wishbone_out[53]
  PIN wishbone_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.530 676.000 471.810 680.000 ;
    END
  END wishbone_out[54]
  PIN wishbone_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.210 676.000 475.490 680.000 ;
    END
  END wishbone_out[55]
  PIN wishbone_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.350 676.000 479.630 680.000 ;
    END
  END wishbone_out[56]
  PIN wishbone_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.030 676.000 483.310 680.000 ;
    END
  END wishbone_out[57]
  PIN wishbone_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.170 676.000 487.450 680.000 ;
    END
  END wishbone_out[58]
  PIN wishbone_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.850 676.000 491.130 680.000 ;
    END
  END wishbone_out[59]
  PIN wishbone_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.790 676.000 279.070 680.000 ;
    END
  END wishbone_out[5]
  PIN wishbone_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.990 676.000 495.270 680.000 ;
    END
  END wishbone_out[60]
  PIN wishbone_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.130 676.000 499.410 680.000 ;
    END
  END wishbone_out[61]
  PIN wishbone_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.810 676.000 503.090 680.000 ;
    END
  END wishbone_out[62]
  PIN wishbone_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.950 676.000 507.230 680.000 ;
    END
  END wishbone_out[63]
  PIN wishbone_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.630 676.000 510.910 680.000 ;
    END
  END wishbone_out[64]
  PIN wishbone_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.770 676.000 515.050 680.000 ;
    END
  END wishbone_out[65]
  PIN wishbone_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.450 676.000 518.730 680.000 ;
    END
  END wishbone_out[66]
  PIN wishbone_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.590 676.000 522.870 680.000 ;
    END
  END wishbone_out[67]
  PIN wishbone_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.270 676.000 526.550 680.000 ;
    END
  END wishbone_out[68]
  PIN wishbone_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.410 676.000 530.690 680.000 ;
    END
  END wishbone_out[69]
  PIN wishbone_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.930 676.000 283.210 680.000 ;
    END
  END wishbone_out[6]
  PIN wishbone_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.090 676.000 534.370 680.000 ;
    END
  END wishbone_out[70]
  PIN wishbone_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.230 676.000 538.510 680.000 ;
    END
  END wishbone_out[71]
  PIN wishbone_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.910 676.000 542.190 680.000 ;
    END
  END wishbone_out[72]
  PIN wishbone_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.050 676.000 546.330 680.000 ;
    END
  END wishbone_out[73]
  PIN wishbone_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.190 676.000 550.470 680.000 ;
    END
  END wishbone_out[74]
  PIN wishbone_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.870 676.000 554.150 680.000 ;
    END
  END wishbone_out[75]
  PIN wishbone_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.010 676.000 558.290 680.000 ;
    END
  END wishbone_out[76]
  PIN wishbone_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.690 676.000 561.970 680.000 ;
    END
  END wishbone_out[77]
  PIN wishbone_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.830 676.000 566.110 680.000 ;
    END
  END wishbone_out[78]
  PIN wishbone_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.510 676.000 569.790 680.000 ;
    END
  END wishbone_out[79]
  PIN wishbone_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.610 676.000 286.890 680.000 ;
    END
  END wishbone_out[7]
  PIN wishbone_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.650 676.000 573.930 680.000 ;
    END
  END wishbone_out[80]
  PIN wishbone_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.330 676.000 577.610 680.000 ;
    END
  END wishbone_out[81]
  PIN wishbone_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.470 676.000 581.750 680.000 ;
    END
  END wishbone_out[82]
  PIN wishbone_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.150 676.000 585.430 680.000 ;
    END
  END wishbone_out[83]
  PIN wishbone_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.290 676.000 589.570 680.000 ;
    END
  END wishbone_out[84]
  PIN wishbone_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.430 676.000 593.710 680.000 ;
    END
  END wishbone_out[85]
  PIN wishbone_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.110 676.000 597.390 680.000 ;
    END
  END wishbone_out[86]
  PIN wishbone_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.250 676.000 601.530 680.000 ;
    END
  END wishbone_out[87]
  PIN wishbone_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.930 676.000 605.210 680.000 ;
    END
  END wishbone_out[88]
  PIN wishbone_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.070 676.000 609.350 680.000 ;
    END
  END wishbone_out[89]
  PIN wishbone_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.750 676.000 291.030 680.000 ;
    END
  END wishbone_out[8]
  PIN wishbone_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.750 676.000 613.030 680.000 ;
    END
  END wishbone_out[90]
  PIN wishbone_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.890 676.000 617.170 680.000 ;
    END
  END wishbone_out[91]
  PIN wishbone_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.570 676.000 620.850 680.000 ;
    END
  END wishbone_out[92]
  PIN wishbone_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.710 676.000 624.990 680.000 ;
    END
  END wishbone_out[93]
  PIN wishbone_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.390 676.000 628.670 680.000 ;
    END
  END wishbone_out[94]
  PIN wishbone_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.530 676.000 632.810 680.000 ;
    END
  END wishbone_out[95]
  PIN wishbone_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.670 676.000 636.950 680.000 ;
    END
  END wishbone_out[96]
  PIN wishbone_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.350 676.000 640.630 680.000 ;
    END
  END wishbone_out[97]
  PIN wishbone_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.490 676.000 644.770 680.000 ;
    END
  END wishbone_out[98]
  PIN wishbone_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.170 676.000 648.450 680.000 ;
    END
  END wishbone_out[99]
  PIN wishbone_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.430 676.000 294.710 680.000 ;
    END
  END wishbone_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 633.540 10.640 635.140 669.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 479.940 10.640 481.540 669.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 326.340 10.640 327.940 669.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 172.740 10.640 174.340 669.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.140 10.640 20.740 669.360 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 556.740 10.640 558.340 669.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 403.140 10.640 404.740 669.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 249.540 10.640 251.140 669.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.940 10.640 97.540 669.360 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 636.840 10.880 638.440 669.120 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 483.240 10.880 484.840 669.120 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 329.640 10.880 331.240 669.120 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 176.040 10.880 177.640 669.120 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.440 10.880 24.040 669.120 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 560.040 10.880 561.640 669.120 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 406.440 10.880 408.040 669.120 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 252.840 10.880 254.440 669.120 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 99.240 10.880 100.840 669.120 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 640.140 10.880 641.740 669.120 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 486.540 10.880 488.140 669.120 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 332.940 10.880 334.540 669.120 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 179.340 10.880 180.940 669.120 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 25.740 10.880 27.340 669.120 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 563.340 10.880 564.940 669.120 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 409.740 10.880 411.340 669.120 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 256.140 10.880 257.740 669.120 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 102.540 10.880 104.140 669.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 643.440 10.880 645.040 669.120 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 489.840 10.880 491.440 669.120 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 336.240 10.880 337.840 669.120 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 182.640 10.880 184.240 669.120 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 29.040 10.880 30.640 669.120 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 566.640 10.880 568.240 669.120 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 413.040 10.880 414.640 669.120 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 259.440 10.880 261.040 669.120 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 105.840 10.880 107.440 669.120 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 3.620 10.795 672.460 669.205 ;
      LAYER met1 ;
        RECT 0.010 0.040 676.070 670.100 ;
      LAYER met2 ;
        RECT 0.590 675.720 3.430 676.000 ;
        RECT 4.270 675.720 7.570 676.000 ;
        RECT 8.410 675.720 11.250 676.000 ;
        RECT 12.090 675.720 15.390 676.000 ;
        RECT 16.230 675.720 19.070 676.000 ;
        RECT 19.910 675.720 23.210 676.000 ;
        RECT 24.050 675.720 26.890 676.000 ;
        RECT 27.730 675.720 31.030 676.000 ;
        RECT 31.870 675.720 34.710 676.000 ;
        RECT 35.550 675.720 38.850 676.000 ;
        RECT 39.690 675.720 42.530 676.000 ;
        RECT 43.370 675.720 46.670 676.000 ;
        RECT 47.510 675.720 50.810 676.000 ;
        RECT 51.650 675.720 54.490 676.000 ;
        RECT 55.330 675.720 58.630 676.000 ;
        RECT 59.470 675.720 62.310 676.000 ;
        RECT 63.150 675.720 66.450 676.000 ;
        RECT 67.290 675.720 70.130 676.000 ;
        RECT 70.970 675.720 74.270 676.000 ;
        RECT 75.110 675.720 77.950 676.000 ;
        RECT 78.790 675.720 82.090 676.000 ;
        RECT 82.930 675.720 85.770 676.000 ;
        RECT 86.610 675.720 89.910 676.000 ;
        RECT 90.750 675.720 94.050 676.000 ;
        RECT 94.890 675.720 97.730 676.000 ;
        RECT 98.570 675.720 101.870 676.000 ;
        RECT 102.710 675.720 105.550 676.000 ;
        RECT 106.390 675.720 109.690 676.000 ;
        RECT 110.530 675.720 113.370 676.000 ;
        RECT 114.210 675.720 117.510 676.000 ;
        RECT 118.350 675.720 121.190 676.000 ;
        RECT 122.030 675.720 125.330 676.000 ;
        RECT 126.170 675.720 129.010 676.000 ;
        RECT 129.850 675.720 133.150 676.000 ;
        RECT 133.990 675.720 137.290 676.000 ;
        RECT 138.130 675.720 140.970 676.000 ;
        RECT 141.810 675.720 145.110 676.000 ;
        RECT 145.950 675.720 148.790 676.000 ;
        RECT 149.630 675.720 152.930 676.000 ;
        RECT 153.770 675.720 156.610 676.000 ;
        RECT 157.450 675.720 160.750 676.000 ;
        RECT 161.590 675.720 164.430 676.000 ;
        RECT 165.270 675.720 168.570 676.000 ;
        RECT 169.410 675.720 172.250 676.000 ;
        RECT 173.090 675.720 176.390 676.000 ;
        RECT 177.230 675.720 180.070 676.000 ;
        RECT 180.910 675.720 184.210 676.000 ;
        RECT 185.050 675.720 188.350 676.000 ;
        RECT 189.190 675.720 192.030 676.000 ;
        RECT 192.870 675.720 196.170 676.000 ;
        RECT 197.010 675.720 199.850 676.000 ;
        RECT 200.690 675.720 203.990 676.000 ;
        RECT 204.830 675.720 207.670 676.000 ;
        RECT 208.510 675.720 211.810 676.000 ;
        RECT 212.650 675.720 215.490 676.000 ;
        RECT 216.330 675.720 219.630 676.000 ;
        RECT 220.470 675.720 223.310 676.000 ;
        RECT 224.150 675.720 227.450 676.000 ;
        RECT 228.290 675.720 231.590 676.000 ;
        RECT 232.430 675.720 235.270 676.000 ;
        RECT 236.110 675.720 239.410 676.000 ;
        RECT 240.250 675.720 243.090 676.000 ;
        RECT 243.930 675.720 247.230 676.000 ;
        RECT 248.070 675.720 250.910 676.000 ;
        RECT 251.750 675.720 255.050 676.000 ;
        RECT 255.890 675.720 258.730 676.000 ;
        RECT 259.570 675.720 262.870 676.000 ;
        RECT 263.710 675.720 266.550 676.000 ;
        RECT 267.390 675.720 270.690 676.000 ;
        RECT 271.530 675.720 274.830 676.000 ;
        RECT 275.670 675.720 278.510 676.000 ;
        RECT 279.350 675.720 282.650 676.000 ;
        RECT 283.490 675.720 286.330 676.000 ;
        RECT 287.170 675.720 290.470 676.000 ;
        RECT 291.310 675.720 294.150 676.000 ;
        RECT 294.990 675.720 298.290 676.000 ;
        RECT 299.130 675.720 301.970 676.000 ;
        RECT 302.810 675.720 306.110 676.000 ;
        RECT 306.950 675.720 309.790 676.000 ;
        RECT 310.630 675.720 313.930 676.000 ;
        RECT 314.770 675.720 318.070 676.000 ;
        RECT 318.910 675.720 321.750 676.000 ;
        RECT 322.590 675.720 325.890 676.000 ;
        RECT 326.730 675.720 329.570 676.000 ;
        RECT 330.410 675.720 333.710 676.000 ;
        RECT 334.550 675.720 337.390 676.000 ;
        RECT 338.230 675.720 341.530 676.000 ;
        RECT 342.370 675.720 345.210 676.000 ;
        RECT 346.050 675.720 349.350 676.000 ;
        RECT 350.190 675.720 353.030 676.000 ;
        RECT 353.870 675.720 357.170 676.000 ;
        RECT 358.010 675.720 360.850 676.000 ;
        RECT 361.690 675.720 364.990 676.000 ;
        RECT 365.830 675.720 369.130 676.000 ;
        RECT 369.970 675.720 372.810 676.000 ;
        RECT 373.650 675.720 376.950 676.000 ;
        RECT 377.790 675.720 380.630 676.000 ;
        RECT 381.470 675.720 384.770 676.000 ;
        RECT 385.610 675.720 388.450 676.000 ;
        RECT 389.290 675.720 392.590 676.000 ;
        RECT 393.430 675.720 396.270 676.000 ;
        RECT 397.110 675.720 400.410 676.000 ;
        RECT 401.250 675.720 404.090 676.000 ;
        RECT 404.930 675.720 408.230 676.000 ;
        RECT 409.070 675.720 412.370 676.000 ;
        RECT 413.210 675.720 416.050 676.000 ;
        RECT 416.890 675.720 420.190 676.000 ;
        RECT 421.030 675.720 423.870 676.000 ;
        RECT 424.710 675.720 428.010 676.000 ;
        RECT 428.850 675.720 431.690 676.000 ;
        RECT 432.530 675.720 435.830 676.000 ;
        RECT 436.670 675.720 439.510 676.000 ;
        RECT 440.350 675.720 443.650 676.000 ;
        RECT 444.490 675.720 447.330 676.000 ;
        RECT 448.170 675.720 451.470 676.000 ;
        RECT 452.310 675.720 455.610 676.000 ;
        RECT 456.450 675.720 459.290 676.000 ;
        RECT 460.130 675.720 463.430 676.000 ;
        RECT 464.270 675.720 467.110 676.000 ;
        RECT 467.950 675.720 471.250 676.000 ;
        RECT 472.090 675.720 474.930 676.000 ;
        RECT 475.770 675.720 479.070 676.000 ;
        RECT 479.910 675.720 482.750 676.000 ;
        RECT 483.590 675.720 486.890 676.000 ;
        RECT 487.730 675.720 490.570 676.000 ;
        RECT 491.410 675.720 494.710 676.000 ;
        RECT 495.550 675.720 498.850 676.000 ;
        RECT 499.690 675.720 502.530 676.000 ;
        RECT 503.370 675.720 506.670 676.000 ;
        RECT 507.510 675.720 510.350 676.000 ;
        RECT 511.190 675.720 514.490 676.000 ;
        RECT 515.330 675.720 518.170 676.000 ;
        RECT 519.010 675.720 522.310 676.000 ;
        RECT 523.150 675.720 525.990 676.000 ;
        RECT 526.830 675.720 530.130 676.000 ;
        RECT 530.970 675.720 533.810 676.000 ;
        RECT 534.650 675.720 537.950 676.000 ;
        RECT 538.790 675.720 541.630 676.000 ;
        RECT 542.470 675.720 545.770 676.000 ;
        RECT 546.610 675.720 549.910 676.000 ;
        RECT 550.750 675.720 553.590 676.000 ;
        RECT 554.430 675.720 557.730 676.000 ;
        RECT 558.570 675.720 561.410 676.000 ;
        RECT 562.250 675.720 565.550 676.000 ;
        RECT 566.390 675.720 569.230 676.000 ;
        RECT 570.070 675.720 573.370 676.000 ;
        RECT 574.210 675.720 577.050 676.000 ;
        RECT 577.890 675.720 581.190 676.000 ;
        RECT 582.030 675.720 584.870 676.000 ;
        RECT 585.710 675.720 589.010 676.000 ;
        RECT 589.850 675.720 593.150 676.000 ;
        RECT 593.990 675.720 596.830 676.000 ;
        RECT 597.670 675.720 600.970 676.000 ;
        RECT 601.810 675.720 604.650 676.000 ;
        RECT 605.490 675.720 608.790 676.000 ;
        RECT 609.630 675.720 612.470 676.000 ;
        RECT 613.310 675.720 616.610 676.000 ;
        RECT 617.450 675.720 620.290 676.000 ;
        RECT 621.130 675.720 624.430 676.000 ;
        RECT 625.270 675.720 628.110 676.000 ;
        RECT 628.950 675.720 632.250 676.000 ;
        RECT 633.090 675.720 636.390 676.000 ;
        RECT 637.230 675.720 640.070 676.000 ;
        RECT 640.910 675.720 644.210 676.000 ;
        RECT 645.050 675.720 647.890 676.000 ;
        RECT 648.730 675.720 652.030 676.000 ;
        RECT 652.870 675.720 655.710 676.000 ;
        RECT 656.550 675.720 659.850 676.000 ;
        RECT 660.690 675.720 663.530 676.000 ;
        RECT 664.370 675.720 667.670 676.000 ;
        RECT 668.510 675.720 671.350 676.000 ;
        RECT 672.190 675.720 675.490 676.000 ;
        RECT 0.030 4.280 676.040 675.720 ;
        RECT 0.590 0.010 3.430 4.280 ;
        RECT 4.270 0.010 7.570 4.280 ;
        RECT 8.410 0.010 11.250 4.280 ;
        RECT 12.090 0.010 15.390 4.280 ;
        RECT 16.230 0.010 19.070 4.280 ;
        RECT 19.910 0.010 23.210 4.280 ;
        RECT 24.050 0.010 26.890 4.280 ;
        RECT 27.730 0.010 31.030 4.280 ;
        RECT 31.870 0.010 34.710 4.280 ;
        RECT 35.550 0.010 38.850 4.280 ;
        RECT 39.690 0.010 42.530 4.280 ;
        RECT 43.370 0.010 46.670 4.280 ;
        RECT 47.510 0.010 50.810 4.280 ;
        RECT 51.650 0.010 54.490 4.280 ;
        RECT 55.330 0.010 58.630 4.280 ;
        RECT 59.470 0.010 62.310 4.280 ;
        RECT 63.150 0.010 66.450 4.280 ;
        RECT 67.290 0.010 70.130 4.280 ;
        RECT 70.970 0.010 74.270 4.280 ;
        RECT 75.110 0.010 77.950 4.280 ;
        RECT 78.790 0.010 82.090 4.280 ;
        RECT 82.930 0.010 85.770 4.280 ;
        RECT 86.610 0.010 89.910 4.280 ;
        RECT 90.750 0.010 94.050 4.280 ;
        RECT 94.890 0.010 97.730 4.280 ;
        RECT 98.570 0.010 101.870 4.280 ;
        RECT 102.710 0.010 105.550 4.280 ;
        RECT 106.390 0.010 109.690 4.280 ;
        RECT 110.530 0.010 113.370 4.280 ;
        RECT 114.210 0.010 117.510 4.280 ;
        RECT 118.350 0.010 121.190 4.280 ;
        RECT 122.030 0.010 125.330 4.280 ;
        RECT 126.170 0.010 129.010 4.280 ;
        RECT 129.850 0.010 133.150 4.280 ;
        RECT 133.990 0.010 137.290 4.280 ;
        RECT 138.130 0.010 140.970 4.280 ;
        RECT 141.810 0.010 145.110 4.280 ;
        RECT 145.950 0.010 148.790 4.280 ;
        RECT 149.630 0.010 152.930 4.280 ;
        RECT 153.770 0.010 156.610 4.280 ;
        RECT 157.450 0.010 160.750 4.280 ;
        RECT 161.590 0.010 164.430 4.280 ;
        RECT 165.270 0.010 168.570 4.280 ;
        RECT 169.410 0.010 172.250 4.280 ;
        RECT 173.090 0.010 176.390 4.280 ;
        RECT 177.230 0.010 180.070 4.280 ;
        RECT 180.910 0.010 184.210 4.280 ;
        RECT 185.050 0.010 188.350 4.280 ;
        RECT 189.190 0.010 192.030 4.280 ;
        RECT 192.870 0.010 196.170 4.280 ;
        RECT 197.010 0.010 199.850 4.280 ;
        RECT 200.690 0.010 203.990 4.280 ;
        RECT 204.830 0.010 207.670 4.280 ;
        RECT 208.510 0.010 211.810 4.280 ;
        RECT 212.650 0.010 215.490 4.280 ;
        RECT 216.330 0.010 219.630 4.280 ;
        RECT 220.470 0.010 223.310 4.280 ;
        RECT 224.150 0.010 227.450 4.280 ;
        RECT 228.290 0.010 231.590 4.280 ;
        RECT 232.430 0.010 235.270 4.280 ;
        RECT 236.110 0.010 239.410 4.280 ;
        RECT 240.250 0.010 243.090 4.280 ;
        RECT 243.930 0.010 247.230 4.280 ;
        RECT 248.070 0.010 250.910 4.280 ;
        RECT 251.750 0.010 255.050 4.280 ;
        RECT 255.890 0.010 258.730 4.280 ;
        RECT 259.570 0.010 262.870 4.280 ;
        RECT 263.710 0.010 266.550 4.280 ;
        RECT 267.390 0.010 270.690 4.280 ;
        RECT 271.530 0.010 274.830 4.280 ;
        RECT 275.670 0.010 278.510 4.280 ;
        RECT 279.350 0.010 282.650 4.280 ;
        RECT 283.490 0.010 286.330 4.280 ;
        RECT 287.170 0.010 290.470 4.280 ;
        RECT 291.310 0.010 294.150 4.280 ;
        RECT 294.990 0.010 298.290 4.280 ;
        RECT 299.130 0.010 301.970 4.280 ;
        RECT 302.810 0.010 306.110 4.280 ;
        RECT 306.950 0.010 309.790 4.280 ;
        RECT 310.630 0.010 313.930 4.280 ;
        RECT 314.770 0.010 318.070 4.280 ;
        RECT 318.910 0.010 321.750 4.280 ;
        RECT 322.590 0.010 325.890 4.280 ;
        RECT 326.730 0.010 329.570 4.280 ;
        RECT 330.410 0.010 333.710 4.280 ;
        RECT 334.550 0.010 337.390 4.280 ;
        RECT 338.230 0.010 341.530 4.280 ;
        RECT 342.370 0.010 345.210 4.280 ;
        RECT 346.050 0.010 349.350 4.280 ;
        RECT 350.190 0.010 353.030 4.280 ;
        RECT 353.870 0.010 357.170 4.280 ;
        RECT 358.010 0.010 360.850 4.280 ;
        RECT 361.690 0.010 364.990 4.280 ;
        RECT 365.830 0.010 369.130 4.280 ;
        RECT 369.970 0.010 372.810 4.280 ;
        RECT 373.650 0.010 376.950 4.280 ;
        RECT 377.790 0.010 380.630 4.280 ;
        RECT 381.470 0.010 384.770 4.280 ;
        RECT 385.610 0.010 388.450 4.280 ;
        RECT 389.290 0.010 392.590 4.280 ;
        RECT 393.430 0.010 396.270 4.280 ;
        RECT 397.110 0.010 400.410 4.280 ;
        RECT 401.250 0.010 404.090 4.280 ;
        RECT 404.930 0.010 408.230 4.280 ;
        RECT 409.070 0.010 412.370 4.280 ;
        RECT 413.210 0.010 416.050 4.280 ;
        RECT 416.890 0.010 420.190 4.280 ;
        RECT 421.030 0.010 423.870 4.280 ;
        RECT 424.710 0.010 428.010 4.280 ;
        RECT 428.850 0.010 431.690 4.280 ;
        RECT 432.530 0.010 435.830 4.280 ;
        RECT 436.670 0.010 439.510 4.280 ;
        RECT 440.350 0.010 443.650 4.280 ;
        RECT 444.490 0.010 447.330 4.280 ;
        RECT 448.170 0.010 451.470 4.280 ;
        RECT 452.310 0.010 455.610 4.280 ;
        RECT 456.450 0.010 459.290 4.280 ;
        RECT 460.130 0.010 463.430 4.280 ;
        RECT 464.270 0.010 467.110 4.280 ;
        RECT 467.950 0.010 471.250 4.280 ;
        RECT 472.090 0.010 474.930 4.280 ;
        RECT 475.770 0.010 479.070 4.280 ;
        RECT 479.910 0.010 482.750 4.280 ;
        RECT 483.590 0.010 486.890 4.280 ;
        RECT 487.730 0.010 490.570 4.280 ;
        RECT 491.410 0.010 494.710 4.280 ;
        RECT 495.550 0.010 498.850 4.280 ;
        RECT 499.690 0.010 502.530 4.280 ;
        RECT 503.370 0.010 506.670 4.280 ;
        RECT 507.510 0.010 510.350 4.280 ;
        RECT 511.190 0.010 514.490 4.280 ;
        RECT 515.330 0.010 518.170 4.280 ;
        RECT 519.010 0.010 522.310 4.280 ;
        RECT 523.150 0.010 525.990 4.280 ;
        RECT 526.830 0.010 530.130 4.280 ;
        RECT 530.970 0.010 533.810 4.280 ;
        RECT 534.650 0.010 537.950 4.280 ;
        RECT 538.790 0.010 541.630 4.280 ;
        RECT 542.470 0.010 545.770 4.280 ;
        RECT 546.610 0.010 549.910 4.280 ;
        RECT 550.750 0.010 553.590 4.280 ;
        RECT 554.430 0.010 557.730 4.280 ;
        RECT 558.570 0.010 561.410 4.280 ;
        RECT 562.250 0.010 565.550 4.280 ;
        RECT 566.390 0.010 569.230 4.280 ;
        RECT 570.070 0.010 573.370 4.280 ;
        RECT 574.210 0.010 577.050 4.280 ;
        RECT 577.890 0.010 581.190 4.280 ;
        RECT 582.030 0.010 584.870 4.280 ;
        RECT 585.710 0.010 589.010 4.280 ;
        RECT 589.850 0.010 593.150 4.280 ;
        RECT 593.990 0.010 596.830 4.280 ;
        RECT 597.670 0.010 600.970 4.280 ;
        RECT 601.810 0.010 604.650 4.280 ;
        RECT 605.490 0.010 608.790 4.280 ;
        RECT 609.630 0.010 612.470 4.280 ;
        RECT 613.310 0.010 616.610 4.280 ;
        RECT 617.450 0.010 620.290 4.280 ;
        RECT 621.130 0.010 624.430 4.280 ;
        RECT 625.270 0.010 628.110 4.280 ;
        RECT 628.950 0.010 632.250 4.280 ;
        RECT 633.090 0.010 636.390 4.280 ;
        RECT 637.230 0.010 640.070 4.280 ;
        RECT 640.910 0.010 644.210 4.280 ;
        RECT 645.050 0.010 647.890 4.280 ;
        RECT 648.730 0.010 652.030 4.280 ;
        RECT 652.870 0.010 655.710 4.280 ;
        RECT 656.550 0.010 659.850 4.280 ;
        RECT 660.690 0.010 663.530 4.280 ;
        RECT 664.370 0.010 667.670 4.280 ;
        RECT 668.510 0.010 671.350 4.280 ;
        RECT 672.190 0.010 675.490 4.280 ;
      LAYER met3 ;
        RECT 0.005 667.440 674.235 670.300 ;
        RECT 0.005 666.040 673.700 667.440 ;
        RECT 0.005 662.000 674.235 666.040 ;
        RECT 0.005 660.600 673.700 662.000 ;
        RECT 0.005 657.240 674.235 660.600 ;
        RECT 0.005 655.840 673.700 657.240 ;
        RECT 0.005 651.800 674.235 655.840 ;
        RECT 0.005 650.400 673.700 651.800 ;
        RECT 0.005 647.040 674.235 650.400 ;
        RECT 0.005 645.640 673.700 647.040 ;
        RECT 0.005 641.600 674.235 645.640 ;
        RECT 0.005 640.200 673.700 641.600 ;
        RECT 0.005 636.840 674.235 640.200 ;
        RECT 0.005 635.440 673.700 636.840 ;
        RECT 0.005 631.400 674.235 635.440 ;
        RECT 0.005 630.000 673.700 631.400 ;
        RECT 0.005 626.640 674.235 630.000 ;
        RECT 0.005 625.240 673.700 626.640 ;
        RECT 0.005 621.200 674.235 625.240 ;
        RECT 0.005 619.800 673.700 621.200 ;
        RECT 0.005 616.440 674.235 619.800 ;
        RECT 0.005 615.040 673.700 616.440 ;
        RECT 0.005 611.000 674.235 615.040 ;
        RECT 0.005 609.600 673.700 611.000 ;
        RECT 0.005 606.240 674.235 609.600 ;
        RECT 0.005 604.840 673.700 606.240 ;
        RECT 0.005 600.800 674.235 604.840 ;
        RECT 0.005 599.400 673.700 600.800 ;
        RECT 0.005 596.040 674.235 599.400 ;
        RECT 0.005 594.640 673.700 596.040 ;
        RECT 0.005 590.600 674.235 594.640 ;
        RECT 0.005 589.200 673.700 590.600 ;
        RECT 0.005 585.840 674.235 589.200 ;
        RECT 0.005 584.440 673.700 585.840 ;
        RECT 0.005 580.400 674.235 584.440 ;
        RECT 0.005 579.000 673.700 580.400 ;
        RECT 0.005 575.640 674.235 579.000 ;
        RECT 0.005 574.240 673.700 575.640 ;
        RECT 0.005 570.200 674.235 574.240 ;
        RECT 0.005 568.800 673.700 570.200 ;
        RECT 0.005 565.440 674.235 568.800 ;
        RECT 0.005 564.040 673.700 565.440 ;
        RECT 0.005 560.000 674.235 564.040 ;
        RECT 0.005 558.600 673.700 560.000 ;
        RECT 0.005 555.240 674.235 558.600 ;
        RECT 0.005 553.840 673.700 555.240 ;
        RECT 0.005 549.800 674.235 553.840 ;
        RECT 0.005 548.400 673.700 549.800 ;
        RECT 0.005 544.360 674.235 548.400 ;
        RECT 0.005 542.960 673.700 544.360 ;
        RECT 0.005 539.600 674.235 542.960 ;
        RECT 0.005 538.200 673.700 539.600 ;
        RECT 0.005 534.160 674.235 538.200 ;
        RECT 0.005 532.760 673.700 534.160 ;
        RECT 0.005 529.400 674.235 532.760 ;
        RECT 0.005 528.000 673.700 529.400 ;
        RECT 0.005 523.960 674.235 528.000 ;
        RECT 0.005 522.560 673.700 523.960 ;
        RECT 0.005 519.200 674.235 522.560 ;
        RECT 0.005 517.800 673.700 519.200 ;
        RECT 0.005 513.760 674.235 517.800 ;
        RECT 0.005 512.360 673.700 513.760 ;
        RECT 0.005 509.000 674.235 512.360 ;
        RECT 0.005 507.600 673.700 509.000 ;
        RECT 0.005 503.560 674.235 507.600 ;
        RECT 0.005 502.160 673.700 503.560 ;
        RECT 0.005 498.800 674.235 502.160 ;
        RECT 0.005 497.400 673.700 498.800 ;
        RECT 0.005 493.360 674.235 497.400 ;
        RECT 0.005 491.960 673.700 493.360 ;
        RECT 0.005 488.600 674.235 491.960 ;
        RECT 0.005 487.200 673.700 488.600 ;
        RECT 0.005 483.160 674.235 487.200 ;
        RECT 0.005 481.760 673.700 483.160 ;
        RECT 0.005 478.400 674.235 481.760 ;
        RECT 0.005 477.000 673.700 478.400 ;
        RECT 0.005 472.960 674.235 477.000 ;
        RECT 0.005 471.560 673.700 472.960 ;
        RECT 0.005 468.200 674.235 471.560 ;
        RECT 0.005 466.800 673.700 468.200 ;
        RECT 0.005 462.760 674.235 466.800 ;
        RECT 0.005 461.360 673.700 462.760 ;
        RECT 0.005 458.000 674.235 461.360 ;
        RECT 0.005 456.600 673.700 458.000 ;
        RECT 0.005 452.560 674.235 456.600 ;
        RECT 0.005 451.160 673.700 452.560 ;
        RECT 0.005 447.800 674.235 451.160 ;
        RECT 0.005 446.400 673.700 447.800 ;
        RECT 0.005 442.360 674.235 446.400 ;
        RECT 0.005 440.960 673.700 442.360 ;
        RECT 0.005 437.600 674.235 440.960 ;
        RECT 0.005 436.200 673.700 437.600 ;
        RECT 0.005 432.160 674.235 436.200 ;
        RECT 0.005 430.760 673.700 432.160 ;
        RECT 0.005 427.400 674.235 430.760 ;
        RECT 0.005 426.000 673.700 427.400 ;
        RECT 0.005 421.960 674.235 426.000 ;
        RECT 0.005 420.560 673.700 421.960 ;
        RECT 0.005 417.200 674.235 420.560 ;
        RECT 0.005 415.800 673.700 417.200 ;
        RECT 0.005 411.760 674.235 415.800 ;
        RECT 0.005 410.360 673.700 411.760 ;
        RECT 0.005 406.320 674.235 410.360 ;
        RECT 0.005 404.920 673.700 406.320 ;
        RECT 0.005 401.560 674.235 404.920 ;
        RECT 0.005 400.160 673.700 401.560 ;
        RECT 0.005 396.120 674.235 400.160 ;
        RECT 0.005 394.720 673.700 396.120 ;
        RECT 0.005 391.360 674.235 394.720 ;
        RECT 0.005 389.960 673.700 391.360 ;
        RECT 0.005 385.920 674.235 389.960 ;
        RECT 0.005 384.520 673.700 385.920 ;
        RECT 0.005 381.160 674.235 384.520 ;
        RECT 0.005 379.760 673.700 381.160 ;
        RECT 0.005 375.720 674.235 379.760 ;
        RECT 0.005 374.320 673.700 375.720 ;
        RECT 0.005 370.960 674.235 374.320 ;
        RECT 0.005 369.560 673.700 370.960 ;
        RECT 0.005 365.520 674.235 369.560 ;
        RECT 0.005 364.120 673.700 365.520 ;
        RECT 0.005 360.760 674.235 364.120 ;
        RECT 0.005 359.360 673.700 360.760 ;
        RECT 0.005 355.320 674.235 359.360 ;
        RECT 0.005 353.920 673.700 355.320 ;
        RECT 0.005 350.560 674.235 353.920 ;
        RECT 0.005 349.160 673.700 350.560 ;
        RECT 0.005 345.120 674.235 349.160 ;
        RECT 0.005 343.720 673.700 345.120 ;
        RECT 0.005 340.360 674.235 343.720 ;
        RECT 0.005 338.960 673.700 340.360 ;
        RECT 0.005 334.920 674.235 338.960 ;
        RECT 0.005 333.520 673.700 334.920 ;
        RECT 0.005 330.160 674.235 333.520 ;
        RECT 0.005 328.760 673.700 330.160 ;
        RECT 0.005 324.720 674.235 328.760 ;
        RECT 0.005 323.320 673.700 324.720 ;
        RECT 0.005 319.960 674.235 323.320 ;
        RECT 0.005 318.560 673.700 319.960 ;
        RECT 0.005 314.520 674.235 318.560 ;
        RECT 0.005 313.120 673.700 314.520 ;
        RECT 0.005 309.760 674.235 313.120 ;
        RECT 0.005 308.360 673.700 309.760 ;
        RECT 0.005 304.320 674.235 308.360 ;
        RECT 0.005 302.920 673.700 304.320 ;
        RECT 0.005 299.560 674.235 302.920 ;
        RECT 0.005 298.160 673.700 299.560 ;
        RECT 0.005 294.120 674.235 298.160 ;
        RECT 0.005 292.720 673.700 294.120 ;
        RECT 0.005 289.360 674.235 292.720 ;
        RECT 0.005 287.960 673.700 289.360 ;
        RECT 0.005 283.920 674.235 287.960 ;
        RECT 0.005 282.520 673.700 283.920 ;
        RECT 0.005 279.160 674.235 282.520 ;
        RECT 0.005 277.760 673.700 279.160 ;
        RECT 0.005 273.720 674.235 277.760 ;
        RECT 0.005 272.320 673.700 273.720 ;
        RECT 0.005 268.280 674.235 272.320 ;
        RECT 0.005 266.880 673.700 268.280 ;
        RECT 0.005 263.520 674.235 266.880 ;
        RECT 0.005 262.120 673.700 263.520 ;
        RECT 0.005 258.080 674.235 262.120 ;
        RECT 0.005 256.680 673.700 258.080 ;
        RECT 0.005 253.320 674.235 256.680 ;
        RECT 0.005 251.920 673.700 253.320 ;
        RECT 0.005 247.880 674.235 251.920 ;
        RECT 0.005 246.480 673.700 247.880 ;
        RECT 0.005 243.120 674.235 246.480 ;
        RECT 0.005 241.720 673.700 243.120 ;
        RECT 0.005 237.680 674.235 241.720 ;
        RECT 0.005 236.280 673.700 237.680 ;
        RECT 0.005 232.920 674.235 236.280 ;
        RECT 0.005 231.520 673.700 232.920 ;
        RECT 0.005 227.480 674.235 231.520 ;
        RECT 0.005 226.080 673.700 227.480 ;
        RECT 0.005 222.720 674.235 226.080 ;
        RECT 0.005 221.320 673.700 222.720 ;
        RECT 0.005 217.280 674.235 221.320 ;
        RECT 0.005 215.880 673.700 217.280 ;
        RECT 0.005 212.520 674.235 215.880 ;
        RECT 0.005 211.120 673.700 212.520 ;
        RECT 0.005 207.080 674.235 211.120 ;
        RECT 0.005 205.680 673.700 207.080 ;
        RECT 0.005 202.320 674.235 205.680 ;
        RECT 0.005 200.920 673.700 202.320 ;
        RECT 0.005 196.880 674.235 200.920 ;
        RECT 0.005 195.480 673.700 196.880 ;
        RECT 0.005 192.120 674.235 195.480 ;
        RECT 0.005 190.720 673.700 192.120 ;
        RECT 0.005 186.680 674.235 190.720 ;
        RECT 0.005 185.280 673.700 186.680 ;
        RECT 0.005 181.920 674.235 185.280 ;
        RECT 0.005 180.520 673.700 181.920 ;
        RECT 0.005 176.480 674.235 180.520 ;
        RECT 0.005 175.080 673.700 176.480 ;
        RECT 0.005 171.720 674.235 175.080 ;
        RECT 0.005 170.320 673.700 171.720 ;
        RECT 0.005 166.280 674.235 170.320 ;
        RECT 0.005 164.880 673.700 166.280 ;
        RECT 0.005 161.520 674.235 164.880 ;
        RECT 0.005 160.120 673.700 161.520 ;
        RECT 0.005 156.080 674.235 160.120 ;
        RECT 0.005 154.680 673.700 156.080 ;
        RECT 0.005 151.320 674.235 154.680 ;
        RECT 0.005 149.920 673.700 151.320 ;
        RECT 0.005 145.880 674.235 149.920 ;
        RECT 0.005 144.480 673.700 145.880 ;
        RECT 0.005 141.120 674.235 144.480 ;
        RECT 0.005 139.720 673.700 141.120 ;
        RECT 0.005 135.680 674.235 139.720 ;
        RECT 0.005 134.280 673.700 135.680 ;
        RECT 0.005 130.240 674.235 134.280 ;
        RECT 0.005 128.840 673.700 130.240 ;
        RECT 0.005 125.480 674.235 128.840 ;
        RECT 0.005 124.080 673.700 125.480 ;
        RECT 0.005 120.040 674.235 124.080 ;
        RECT 0.005 118.640 673.700 120.040 ;
        RECT 0.005 115.280 674.235 118.640 ;
        RECT 0.005 113.880 673.700 115.280 ;
        RECT 0.005 109.840 674.235 113.880 ;
        RECT 0.005 108.440 673.700 109.840 ;
        RECT 0.005 105.080 674.235 108.440 ;
        RECT 0.005 103.680 673.700 105.080 ;
        RECT 0.005 99.640 674.235 103.680 ;
        RECT 0.005 98.240 673.700 99.640 ;
        RECT 0.005 94.880 674.235 98.240 ;
        RECT 0.005 93.480 673.700 94.880 ;
        RECT 0.005 89.440 674.235 93.480 ;
        RECT 0.005 88.040 673.700 89.440 ;
        RECT 0.005 84.680 674.235 88.040 ;
        RECT 0.005 83.280 673.700 84.680 ;
        RECT 0.005 79.240 674.235 83.280 ;
        RECT 0.005 77.840 673.700 79.240 ;
        RECT 0.005 74.480 674.235 77.840 ;
        RECT 0.005 73.080 673.700 74.480 ;
        RECT 0.005 69.040 674.235 73.080 ;
        RECT 0.005 67.640 673.700 69.040 ;
        RECT 0.005 64.280 674.235 67.640 ;
        RECT 0.005 62.880 673.700 64.280 ;
        RECT 0.005 58.840 674.235 62.880 ;
        RECT 0.005 57.440 673.700 58.840 ;
        RECT 0.005 54.080 674.235 57.440 ;
        RECT 0.005 52.680 673.700 54.080 ;
        RECT 0.005 48.640 674.235 52.680 ;
        RECT 0.005 47.240 673.700 48.640 ;
        RECT 0.005 43.880 674.235 47.240 ;
        RECT 0.005 42.480 673.700 43.880 ;
        RECT 0.005 38.440 674.235 42.480 ;
        RECT 0.005 37.040 673.700 38.440 ;
        RECT 0.005 33.680 674.235 37.040 ;
        RECT 0.005 32.280 673.700 33.680 ;
        RECT 0.005 28.240 674.235 32.280 ;
        RECT 0.005 26.840 673.700 28.240 ;
        RECT 0.005 23.480 674.235 26.840 ;
        RECT 0.005 22.080 673.700 23.480 ;
        RECT 0.005 18.040 674.235 22.080 ;
        RECT 0.005 16.640 673.700 18.040 ;
        RECT 0.005 13.280 674.235 16.640 ;
        RECT 0.005 11.880 673.700 13.280 ;
        RECT 0.005 7.840 674.235 11.880 ;
        RECT 0.005 6.440 673.700 7.840 ;
        RECT 0.005 3.080 674.235 6.440 ;
        RECT 0.005 1.680 673.700 3.080 ;
        RECT 0.005 0.175 674.235 1.680 ;
      LAYER met4 ;
        RECT 14.035 669.760 666.645 670.305 ;
        RECT 14.035 14.455 18.740 669.760 ;
        RECT 21.140 669.520 95.540 669.760 ;
        RECT 21.140 14.455 22.040 669.520 ;
        RECT 24.440 14.455 25.340 669.520 ;
        RECT 27.740 14.455 28.640 669.520 ;
        RECT 31.040 14.455 95.540 669.520 ;
        RECT 97.940 669.520 172.340 669.760 ;
        RECT 97.940 14.455 98.840 669.520 ;
        RECT 101.240 14.455 102.140 669.520 ;
        RECT 104.540 14.455 105.440 669.520 ;
        RECT 107.840 14.455 172.340 669.520 ;
        RECT 174.740 669.520 249.140 669.760 ;
        RECT 174.740 14.455 175.640 669.520 ;
        RECT 178.040 14.455 178.940 669.520 ;
        RECT 181.340 14.455 182.240 669.520 ;
        RECT 184.640 14.455 249.140 669.520 ;
        RECT 251.540 669.520 325.940 669.760 ;
        RECT 251.540 14.455 252.440 669.520 ;
        RECT 254.840 14.455 255.740 669.520 ;
        RECT 258.140 14.455 259.040 669.520 ;
        RECT 261.440 14.455 325.940 669.520 ;
        RECT 328.340 669.520 402.740 669.760 ;
        RECT 328.340 14.455 329.240 669.520 ;
        RECT 331.640 14.455 332.540 669.520 ;
        RECT 334.940 14.455 335.840 669.520 ;
        RECT 338.240 14.455 402.740 669.520 ;
        RECT 405.140 669.520 479.540 669.760 ;
        RECT 405.140 14.455 406.040 669.520 ;
        RECT 408.440 14.455 409.340 669.520 ;
        RECT 411.740 14.455 412.640 669.520 ;
        RECT 415.040 14.455 479.540 669.520 ;
        RECT 481.940 669.520 556.340 669.760 ;
        RECT 481.940 14.455 482.840 669.520 ;
        RECT 485.240 14.455 486.140 669.520 ;
        RECT 488.540 14.455 489.440 669.520 ;
        RECT 491.840 14.455 556.340 669.520 ;
        RECT 558.740 669.520 633.140 669.760 ;
        RECT 558.740 14.455 559.640 669.520 ;
        RECT 562.040 14.455 562.940 669.520 ;
        RECT 565.340 14.455 566.240 669.520 ;
        RECT 568.640 14.455 633.140 669.520 ;
        RECT 635.540 669.520 666.645 669.760 ;
        RECT 635.540 14.455 636.440 669.520 ;
        RECT 638.840 14.455 639.740 669.520 ;
        RECT 642.140 14.455 643.040 669.520 ;
        RECT 645.440 14.455 666.645 669.520 ;
  END
END icache
END LIBRARY

