magic
tech sky130A
magscale 1 2
timestamp 1610962084
<< obsli1 >>
rect 724 2159 134492 133841
<< obsm1 >>
rect 2 8 135214 134020
<< metal2 >>
rect 6 135200 62 136000
rect 742 135200 798 136000
rect 1570 135200 1626 136000
rect 2306 135200 2362 136000
rect 3134 135200 3190 136000
rect 3870 135200 3926 136000
rect 4698 135200 4754 136000
rect 5434 135200 5490 136000
rect 6262 135200 6318 136000
rect 6998 135200 7054 136000
rect 7826 135200 7882 136000
rect 8562 135200 8618 136000
rect 9390 135200 9446 136000
rect 10218 135200 10274 136000
rect 10954 135200 11010 136000
rect 11782 135200 11838 136000
rect 12518 135200 12574 136000
rect 13346 135200 13402 136000
rect 14082 135200 14138 136000
rect 14910 135200 14966 136000
rect 15646 135200 15702 136000
rect 16474 135200 16530 136000
rect 17210 135200 17266 136000
rect 18038 135200 18094 136000
rect 18866 135200 18922 136000
rect 19602 135200 19658 136000
rect 20430 135200 20486 136000
rect 21166 135200 21222 136000
rect 21994 135200 22050 136000
rect 22730 135200 22786 136000
rect 23558 135200 23614 136000
rect 24294 135200 24350 136000
rect 25122 135200 25178 136000
rect 25858 135200 25914 136000
rect 26686 135200 26742 136000
rect 27514 135200 27570 136000
rect 28250 135200 28306 136000
rect 29078 135200 29134 136000
rect 29814 135200 29870 136000
rect 30642 135200 30698 136000
rect 31378 135200 31434 136000
rect 32206 135200 32262 136000
rect 32942 135200 32998 136000
rect 33770 135200 33826 136000
rect 34506 135200 34562 136000
rect 35334 135200 35390 136000
rect 36070 135200 36126 136000
rect 36898 135200 36954 136000
rect 37726 135200 37782 136000
rect 38462 135200 38518 136000
rect 39290 135200 39346 136000
rect 40026 135200 40082 136000
rect 40854 135200 40910 136000
rect 41590 135200 41646 136000
rect 42418 135200 42474 136000
rect 43154 135200 43210 136000
rect 43982 135200 44038 136000
rect 44718 135200 44774 136000
rect 45546 135200 45602 136000
rect 46374 135200 46430 136000
rect 47110 135200 47166 136000
rect 47938 135200 47994 136000
rect 48674 135200 48730 136000
rect 49502 135200 49558 136000
rect 50238 135200 50294 136000
rect 51066 135200 51122 136000
rect 51802 135200 51858 136000
rect 52630 135200 52686 136000
rect 53366 135200 53422 136000
rect 54194 135200 54250 136000
rect 55022 135200 55078 136000
rect 55758 135200 55814 136000
rect 56586 135200 56642 136000
rect 57322 135200 57378 136000
rect 58150 135200 58206 136000
rect 58886 135200 58942 136000
rect 59714 135200 59770 136000
rect 60450 135200 60506 136000
rect 61278 135200 61334 136000
rect 62014 135200 62070 136000
rect 62842 135200 62898 136000
rect 63670 135200 63726 136000
rect 64406 135200 64462 136000
rect 65234 135200 65290 136000
rect 65970 135200 66026 136000
rect 66798 135200 66854 136000
rect 67534 135200 67590 136000
rect 68362 135200 68418 136000
rect 69098 135200 69154 136000
rect 69926 135200 69982 136000
rect 70662 135200 70718 136000
rect 71490 135200 71546 136000
rect 72226 135200 72282 136000
rect 73054 135200 73110 136000
rect 73882 135200 73938 136000
rect 74618 135200 74674 136000
rect 75446 135200 75502 136000
rect 76182 135200 76238 136000
rect 77010 135200 77066 136000
rect 77746 135200 77802 136000
rect 78574 135200 78630 136000
rect 79310 135200 79366 136000
rect 80138 135200 80194 136000
rect 80874 135200 80930 136000
rect 81702 135200 81758 136000
rect 82530 135200 82586 136000
rect 83266 135200 83322 136000
rect 84094 135200 84150 136000
rect 84830 135200 84886 136000
rect 85658 135200 85714 136000
rect 86394 135200 86450 136000
rect 87222 135200 87278 136000
rect 87958 135200 88014 136000
rect 88786 135200 88842 136000
rect 89522 135200 89578 136000
rect 90350 135200 90406 136000
rect 91178 135200 91234 136000
rect 91914 135200 91970 136000
rect 92742 135200 92798 136000
rect 93478 135200 93534 136000
rect 94306 135200 94362 136000
rect 95042 135200 95098 136000
rect 95870 135200 95926 136000
rect 96606 135200 96662 136000
rect 97434 135200 97490 136000
rect 98170 135200 98226 136000
rect 98998 135200 99054 136000
rect 99826 135200 99882 136000
rect 100562 135200 100618 136000
rect 101390 135200 101446 136000
rect 102126 135200 102182 136000
rect 102954 135200 103010 136000
rect 103690 135200 103746 136000
rect 104518 135200 104574 136000
rect 105254 135200 105310 136000
rect 106082 135200 106138 136000
rect 106818 135200 106874 136000
rect 107646 135200 107702 136000
rect 108382 135200 108438 136000
rect 109210 135200 109266 136000
rect 110038 135200 110094 136000
rect 110774 135200 110830 136000
rect 111602 135200 111658 136000
rect 112338 135200 112394 136000
rect 113166 135200 113222 136000
rect 113902 135200 113958 136000
rect 114730 135200 114786 136000
rect 115466 135200 115522 136000
rect 116294 135200 116350 136000
rect 117030 135200 117086 136000
rect 117858 135200 117914 136000
rect 118686 135200 118742 136000
rect 119422 135200 119478 136000
rect 120250 135200 120306 136000
rect 120986 135200 121042 136000
rect 121814 135200 121870 136000
rect 122550 135200 122606 136000
rect 123378 135200 123434 136000
rect 124114 135200 124170 136000
rect 124942 135200 124998 136000
rect 125678 135200 125734 136000
rect 126506 135200 126562 136000
rect 127334 135200 127390 136000
rect 128070 135200 128126 136000
rect 128898 135200 128954 136000
rect 129634 135200 129690 136000
rect 130462 135200 130518 136000
rect 131198 135200 131254 136000
rect 132026 135200 132082 136000
rect 132762 135200 132818 136000
rect 133590 135200 133646 136000
rect 134326 135200 134382 136000
rect 135154 135200 135210 136000
rect 6 0 62 800
rect 742 0 798 800
rect 1570 0 1626 800
rect 2306 0 2362 800
rect 3134 0 3190 800
rect 3870 0 3926 800
rect 4698 0 4754 800
rect 5434 0 5490 800
rect 6262 0 6318 800
rect 6998 0 7054 800
rect 7826 0 7882 800
rect 8562 0 8618 800
rect 9390 0 9446 800
rect 10218 0 10274 800
rect 10954 0 11010 800
rect 11782 0 11838 800
rect 12518 0 12574 800
rect 13346 0 13402 800
rect 14082 0 14138 800
rect 14910 0 14966 800
rect 15646 0 15702 800
rect 16474 0 16530 800
rect 17210 0 17266 800
rect 18038 0 18094 800
rect 18866 0 18922 800
rect 19602 0 19658 800
rect 20430 0 20486 800
rect 21166 0 21222 800
rect 21994 0 22050 800
rect 22730 0 22786 800
rect 23558 0 23614 800
rect 24294 0 24350 800
rect 25122 0 25178 800
rect 25858 0 25914 800
rect 26686 0 26742 800
rect 27514 0 27570 800
rect 28250 0 28306 800
rect 29078 0 29134 800
rect 29814 0 29870 800
rect 30642 0 30698 800
rect 31378 0 31434 800
rect 32206 0 32262 800
rect 32942 0 32998 800
rect 33770 0 33826 800
rect 34506 0 34562 800
rect 35334 0 35390 800
rect 36070 0 36126 800
rect 36898 0 36954 800
rect 37726 0 37782 800
rect 38462 0 38518 800
rect 39290 0 39346 800
rect 40026 0 40082 800
rect 40854 0 40910 800
rect 41590 0 41646 800
rect 42418 0 42474 800
rect 43154 0 43210 800
rect 43982 0 44038 800
rect 44718 0 44774 800
rect 45546 0 45602 800
rect 46374 0 46430 800
rect 47110 0 47166 800
rect 47938 0 47994 800
rect 48674 0 48730 800
rect 49502 0 49558 800
rect 50238 0 50294 800
rect 51066 0 51122 800
rect 51802 0 51858 800
rect 52630 0 52686 800
rect 53366 0 53422 800
rect 54194 0 54250 800
rect 55022 0 55078 800
rect 55758 0 55814 800
rect 56586 0 56642 800
rect 57322 0 57378 800
rect 58150 0 58206 800
rect 58886 0 58942 800
rect 59714 0 59770 800
rect 60450 0 60506 800
rect 61278 0 61334 800
rect 62014 0 62070 800
rect 62842 0 62898 800
rect 63670 0 63726 800
rect 64406 0 64462 800
rect 65234 0 65290 800
rect 65970 0 66026 800
rect 66798 0 66854 800
rect 67534 0 67590 800
rect 68362 0 68418 800
rect 69098 0 69154 800
rect 69926 0 69982 800
rect 70662 0 70718 800
rect 71490 0 71546 800
rect 72226 0 72282 800
rect 73054 0 73110 800
rect 73882 0 73938 800
rect 74618 0 74674 800
rect 75446 0 75502 800
rect 76182 0 76238 800
rect 77010 0 77066 800
rect 77746 0 77802 800
rect 78574 0 78630 800
rect 79310 0 79366 800
rect 80138 0 80194 800
rect 80874 0 80930 800
rect 81702 0 81758 800
rect 82530 0 82586 800
rect 83266 0 83322 800
rect 84094 0 84150 800
rect 84830 0 84886 800
rect 85658 0 85714 800
rect 86394 0 86450 800
rect 87222 0 87278 800
rect 87958 0 88014 800
rect 88786 0 88842 800
rect 89522 0 89578 800
rect 90350 0 90406 800
rect 91178 0 91234 800
rect 91914 0 91970 800
rect 92742 0 92798 800
rect 93478 0 93534 800
rect 94306 0 94362 800
rect 95042 0 95098 800
rect 95870 0 95926 800
rect 96606 0 96662 800
rect 97434 0 97490 800
rect 98170 0 98226 800
rect 98998 0 99054 800
rect 99826 0 99882 800
rect 100562 0 100618 800
rect 101390 0 101446 800
rect 102126 0 102182 800
rect 102954 0 103010 800
rect 103690 0 103746 800
rect 104518 0 104574 800
rect 105254 0 105310 800
rect 106082 0 106138 800
rect 106818 0 106874 800
rect 107646 0 107702 800
rect 108382 0 108438 800
rect 109210 0 109266 800
rect 110038 0 110094 800
rect 110774 0 110830 800
rect 111602 0 111658 800
rect 112338 0 112394 800
rect 113166 0 113222 800
rect 113902 0 113958 800
rect 114730 0 114786 800
rect 115466 0 115522 800
rect 116294 0 116350 800
rect 117030 0 117086 800
rect 117858 0 117914 800
rect 118686 0 118742 800
rect 119422 0 119478 800
rect 120250 0 120306 800
rect 120986 0 121042 800
rect 121814 0 121870 800
rect 122550 0 122606 800
rect 123378 0 123434 800
rect 124114 0 124170 800
rect 124942 0 124998 800
rect 125678 0 125734 800
rect 126506 0 126562 800
rect 127334 0 127390 800
rect 128070 0 128126 800
rect 128898 0 128954 800
rect 129634 0 129690 800
rect 130462 0 130518 800
rect 131198 0 131254 800
rect 132026 0 132082 800
rect 132762 0 132818 800
rect 133590 0 133646 800
rect 134326 0 134382 800
rect 135154 0 135210 800
<< obsm2 >>
rect 118 135144 686 135200
rect 854 135144 1514 135200
rect 1682 135144 2250 135200
rect 2418 135144 3078 135200
rect 3246 135144 3814 135200
rect 3982 135144 4642 135200
rect 4810 135144 5378 135200
rect 5546 135144 6206 135200
rect 6374 135144 6942 135200
rect 7110 135144 7770 135200
rect 7938 135144 8506 135200
rect 8674 135144 9334 135200
rect 9502 135144 10162 135200
rect 10330 135144 10898 135200
rect 11066 135144 11726 135200
rect 11894 135144 12462 135200
rect 12630 135144 13290 135200
rect 13458 135144 14026 135200
rect 14194 135144 14854 135200
rect 15022 135144 15590 135200
rect 15758 135144 16418 135200
rect 16586 135144 17154 135200
rect 17322 135144 17982 135200
rect 18150 135144 18810 135200
rect 18978 135144 19546 135200
rect 19714 135144 20374 135200
rect 20542 135144 21110 135200
rect 21278 135144 21938 135200
rect 22106 135144 22674 135200
rect 22842 135144 23502 135200
rect 23670 135144 24238 135200
rect 24406 135144 25066 135200
rect 25234 135144 25802 135200
rect 25970 135144 26630 135200
rect 26798 135144 27458 135200
rect 27626 135144 28194 135200
rect 28362 135144 29022 135200
rect 29190 135144 29758 135200
rect 29926 135144 30586 135200
rect 30754 135144 31322 135200
rect 31490 135144 32150 135200
rect 32318 135144 32886 135200
rect 33054 135144 33714 135200
rect 33882 135144 34450 135200
rect 34618 135144 35278 135200
rect 35446 135144 36014 135200
rect 36182 135144 36842 135200
rect 37010 135144 37670 135200
rect 37838 135144 38406 135200
rect 38574 135144 39234 135200
rect 39402 135144 39970 135200
rect 40138 135144 40798 135200
rect 40966 135144 41534 135200
rect 41702 135144 42362 135200
rect 42530 135144 43098 135200
rect 43266 135144 43926 135200
rect 44094 135144 44662 135200
rect 44830 135144 45490 135200
rect 45658 135144 46318 135200
rect 46486 135144 47054 135200
rect 47222 135144 47882 135200
rect 48050 135144 48618 135200
rect 48786 135144 49446 135200
rect 49614 135144 50182 135200
rect 50350 135144 51010 135200
rect 51178 135144 51746 135200
rect 51914 135144 52574 135200
rect 52742 135144 53310 135200
rect 53478 135144 54138 135200
rect 54306 135144 54966 135200
rect 55134 135144 55702 135200
rect 55870 135144 56530 135200
rect 56698 135144 57266 135200
rect 57434 135144 58094 135200
rect 58262 135144 58830 135200
rect 58998 135144 59658 135200
rect 59826 135144 60394 135200
rect 60562 135144 61222 135200
rect 61390 135144 61958 135200
rect 62126 135144 62786 135200
rect 62954 135144 63614 135200
rect 63782 135144 64350 135200
rect 64518 135144 65178 135200
rect 65346 135144 65914 135200
rect 66082 135144 66742 135200
rect 66910 135144 67478 135200
rect 67646 135144 68306 135200
rect 68474 135144 69042 135200
rect 69210 135144 69870 135200
rect 70038 135144 70606 135200
rect 70774 135144 71434 135200
rect 71602 135144 72170 135200
rect 72338 135144 72998 135200
rect 73166 135144 73826 135200
rect 73994 135144 74562 135200
rect 74730 135144 75390 135200
rect 75558 135144 76126 135200
rect 76294 135144 76954 135200
rect 77122 135144 77690 135200
rect 77858 135144 78518 135200
rect 78686 135144 79254 135200
rect 79422 135144 80082 135200
rect 80250 135144 80818 135200
rect 80986 135144 81646 135200
rect 81814 135144 82474 135200
rect 82642 135144 83210 135200
rect 83378 135144 84038 135200
rect 84206 135144 84774 135200
rect 84942 135144 85602 135200
rect 85770 135144 86338 135200
rect 86506 135144 87166 135200
rect 87334 135144 87902 135200
rect 88070 135144 88730 135200
rect 88898 135144 89466 135200
rect 89634 135144 90294 135200
rect 90462 135144 91122 135200
rect 91290 135144 91858 135200
rect 92026 135144 92686 135200
rect 92854 135144 93422 135200
rect 93590 135144 94250 135200
rect 94418 135144 94986 135200
rect 95154 135144 95814 135200
rect 95982 135144 96550 135200
rect 96718 135144 97378 135200
rect 97546 135144 98114 135200
rect 98282 135144 98942 135200
rect 99110 135144 99770 135200
rect 99938 135144 100506 135200
rect 100674 135144 101334 135200
rect 101502 135144 102070 135200
rect 102238 135144 102898 135200
rect 103066 135144 103634 135200
rect 103802 135144 104462 135200
rect 104630 135144 105198 135200
rect 105366 135144 106026 135200
rect 106194 135144 106762 135200
rect 106930 135144 107590 135200
rect 107758 135144 108326 135200
rect 108494 135144 109154 135200
rect 109322 135144 109982 135200
rect 110150 135144 110718 135200
rect 110886 135144 111546 135200
rect 111714 135144 112282 135200
rect 112450 135144 113110 135200
rect 113278 135144 113846 135200
rect 114014 135144 114674 135200
rect 114842 135144 115410 135200
rect 115578 135144 116238 135200
rect 116406 135144 116974 135200
rect 117142 135144 117802 135200
rect 117970 135144 118630 135200
rect 118798 135144 119366 135200
rect 119534 135144 120194 135200
rect 120362 135144 120930 135200
rect 121098 135144 121758 135200
rect 121926 135144 122494 135200
rect 122662 135144 123322 135200
rect 123490 135144 124058 135200
rect 124226 135144 124886 135200
rect 125054 135144 125622 135200
rect 125790 135144 126450 135200
rect 126618 135144 127278 135200
rect 127446 135144 128014 135200
rect 128182 135144 128842 135200
rect 129010 135144 129578 135200
rect 129746 135144 130406 135200
rect 130574 135144 131142 135200
rect 131310 135144 131970 135200
rect 132138 135144 132706 135200
rect 132874 135144 133534 135200
rect 133702 135144 134270 135200
rect 134438 135144 135098 135200
rect 6 856 135208 135144
rect 118 2 686 856
rect 854 2 1514 856
rect 1682 2 2250 856
rect 2418 2 3078 856
rect 3246 2 3814 856
rect 3982 2 4642 856
rect 4810 2 5378 856
rect 5546 2 6206 856
rect 6374 2 6942 856
rect 7110 2 7770 856
rect 7938 2 8506 856
rect 8674 2 9334 856
rect 9502 2 10162 856
rect 10330 2 10898 856
rect 11066 2 11726 856
rect 11894 2 12462 856
rect 12630 2 13290 856
rect 13458 2 14026 856
rect 14194 2 14854 856
rect 15022 2 15590 856
rect 15758 2 16418 856
rect 16586 2 17154 856
rect 17322 2 17982 856
rect 18150 2 18810 856
rect 18978 2 19546 856
rect 19714 2 20374 856
rect 20542 2 21110 856
rect 21278 2 21938 856
rect 22106 2 22674 856
rect 22842 2 23502 856
rect 23670 2 24238 856
rect 24406 2 25066 856
rect 25234 2 25802 856
rect 25970 2 26630 856
rect 26798 2 27458 856
rect 27626 2 28194 856
rect 28362 2 29022 856
rect 29190 2 29758 856
rect 29926 2 30586 856
rect 30754 2 31322 856
rect 31490 2 32150 856
rect 32318 2 32886 856
rect 33054 2 33714 856
rect 33882 2 34450 856
rect 34618 2 35278 856
rect 35446 2 36014 856
rect 36182 2 36842 856
rect 37010 2 37670 856
rect 37838 2 38406 856
rect 38574 2 39234 856
rect 39402 2 39970 856
rect 40138 2 40798 856
rect 40966 2 41534 856
rect 41702 2 42362 856
rect 42530 2 43098 856
rect 43266 2 43926 856
rect 44094 2 44662 856
rect 44830 2 45490 856
rect 45658 2 46318 856
rect 46486 2 47054 856
rect 47222 2 47882 856
rect 48050 2 48618 856
rect 48786 2 49446 856
rect 49614 2 50182 856
rect 50350 2 51010 856
rect 51178 2 51746 856
rect 51914 2 52574 856
rect 52742 2 53310 856
rect 53478 2 54138 856
rect 54306 2 54966 856
rect 55134 2 55702 856
rect 55870 2 56530 856
rect 56698 2 57266 856
rect 57434 2 58094 856
rect 58262 2 58830 856
rect 58998 2 59658 856
rect 59826 2 60394 856
rect 60562 2 61222 856
rect 61390 2 61958 856
rect 62126 2 62786 856
rect 62954 2 63614 856
rect 63782 2 64350 856
rect 64518 2 65178 856
rect 65346 2 65914 856
rect 66082 2 66742 856
rect 66910 2 67478 856
rect 67646 2 68306 856
rect 68474 2 69042 856
rect 69210 2 69870 856
rect 70038 2 70606 856
rect 70774 2 71434 856
rect 71602 2 72170 856
rect 72338 2 72998 856
rect 73166 2 73826 856
rect 73994 2 74562 856
rect 74730 2 75390 856
rect 75558 2 76126 856
rect 76294 2 76954 856
rect 77122 2 77690 856
rect 77858 2 78518 856
rect 78686 2 79254 856
rect 79422 2 80082 856
rect 80250 2 80818 856
rect 80986 2 81646 856
rect 81814 2 82474 856
rect 82642 2 83210 856
rect 83378 2 84038 856
rect 84206 2 84774 856
rect 84942 2 85602 856
rect 85770 2 86338 856
rect 86506 2 87166 856
rect 87334 2 87902 856
rect 88070 2 88730 856
rect 88898 2 89466 856
rect 89634 2 90294 856
rect 90462 2 91122 856
rect 91290 2 91858 856
rect 92026 2 92686 856
rect 92854 2 93422 856
rect 93590 2 94250 856
rect 94418 2 94986 856
rect 95154 2 95814 856
rect 95982 2 96550 856
rect 96718 2 97378 856
rect 97546 2 98114 856
rect 98282 2 98942 856
rect 99110 2 99770 856
rect 99938 2 100506 856
rect 100674 2 101334 856
rect 101502 2 102070 856
rect 102238 2 102898 856
rect 103066 2 103634 856
rect 103802 2 104462 856
rect 104630 2 105198 856
rect 105366 2 106026 856
rect 106194 2 106762 856
rect 106930 2 107590 856
rect 107758 2 108326 856
rect 108494 2 109154 856
rect 109322 2 109982 856
rect 110150 2 110718 856
rect 110886 2 111546 856
rect 111714 2 112282 856
rect 112450 2 113110 856
rect 113278 2 113846 856
rect 114014 2 114674 856
rect 114842 2 115410 856
rect 115578 2 116238 856
rect 116406 2 116974 856
rect 117142 2 117802 856
rect 117970 2 118630 856
rect 118798 2 119366 856
rect 119534 2 120194 856
rect 120362 2 120930 856
rect 121098 2 121758 856
rect 121926 2 122494 856
rect 122662 2 123322 856
rect 123490 2 124058 856
rect 124226 2 124886 856
rect 125054 2 125622 856
rect 125790 2 126450 856
rect 126618 2 127278 856
rect 127446 2 128014 856
rect 128182 2 128842 856
rect 129010 2 129578 856
rect 129746 2 130406 856
rect 130574 2 131142 856
rect 131310 2 131970 856
rect 132138 2 132706 856
rect 132874 2 133534 856
rect 133702 2 134270 856
rect 134438 2 135098 856
<< metal3 >>
rect 134820 135328 135620 135448
rect 134820 134240 135620 134360
rect 134820 133288 135620 133408
rect 134820 132200 135620 132320
rect 134820 131248 135620 131368
rect 134820 130160 135620 130280
rect 134820 129208 135620 129328
rect 134820 128120 135620 128240
rect 134820 127168 135620 127288
rect 134820 126080 135620 126200
rect 134820 125128 135620 125248
rect 134820 124040 135620 124160
rect 134820 123088 135620 123208
rect 134820 122000 135620 122120
rect 134820 121048 135620 121168
rect 134820 119960 135620 120080
rect 134820 119008 135620 119128
rect 134820 117920 135620 118040
rect 134820 116968 135620 117088
rect 134820 115880 135620 116000
rect 134820 114928 135620 115048
rect 134820 113840 135620 113960
rect 134820 112888 135620 113008
rect 134820 111800 135620 111920
rect 134820 110848 135620 110968
rect 134820 109760 135620 109880
rect 134820 108672 135620 108792
rect 134820 107720 135620 107840
rect 134820 106632 135620 106752
rect 134820 105680 135620 105800
rect 134820 104592 135620 104712
rect 134820 103640 135620 103760
rect 134820 102552 135620 102672
rect 134820 101600 135620 101720
rect 134820 100512 135620 100632
rect 134820 99560 135620 99680
rect 134820 98472 135620 98592
rect 134820 97520 135620 97640
rect 134820 96432 135620 96552
rect 134820 95480 135620 95600
rect 134820 94392 135620 94512
rect 134820 93440 135620 93560
rect 134820 92352 135620 92472
rect 134820 91400 135620 91520
rect 134820 90312 135620 90432
rect 134820 89360 135620 89480
rect 134820 88272 135620 88392
rect 134820 87320 135620 87440
rect 134820 86232 135620 86352
rect 134820 85280 135620 85400
rect 134820 84192 135620 84312
rect 134820 83240 135620 83360
rect 134820 82152 135620 82272
rect 134820 81064 135620 81184
rect 134820 80112 135620 80232
rect 134820 79024 135620 79144
rect 134820 78072 135620 78192
rect 134820 76984 135620 77104
rect 134820 76032 135620 76152
rect 134820 74944 135620 75064
rect 134820 73992 135620 74112
rect 134820 72904 135620 73024
rect 134820 71952 135620 72072
rect 134820 70864 135620 70984
rect 134820 69912 135620 70032
rect 134820 68824 135620 68944
rect 134820 67872 135620 67992
rect 134820 66784 135620 66904
rect 134820 65832 135620 65952
rect 134820 64744 135620 64864
rect 134820 63792 135620 63912
rect 134820 62704 135620 62824
rect 134820 61752 135620 61872
rect 134820 60664 135620 60784
rect 134820 59712 135620 59832
rect 134820 58624 135620 58744
rect 134820 57672 135620 57792
rect 134820 56584 135620 56704
rect 134820 55632 135620 55752
rect 134820 54544 135620 54664
rect 134820 53456 135620 53576
rect 134820 52504 135620 52624
rect 134820 51416 135620 51536
rect 134820 50464 135620 50584
rect 134820 49376 135620 49496
rect 134820 48424 135620 48544
rect 134820 47336 135620 47456
rect 134820 46384 135620 46504
rect 134820 45296 135620 45416
rect 134820 44344 135620 44464
rect 134820 43256 135620 43376
rect 134820 42304 135620 42424
rect 134820 41216 135620 41336
rect 134820 40264 135620 40384
rect 134820 39176 135620 39296
rect 134820 38224 135620 38344
rect 134820 37136 135620 37256
rect 134820 36184 135620 36304
rect 134820 35096 135620 35216
rect 134820 34144 135620 34264
rect 134820 33056 135620 33176
rect 134820 32104 135620 32224
rect 134820 31016 135620 31136
rect 134820 30064 135620 30184
rect 134820 28976 135620 29096
rect 134820 28024 135620 28144
rect 134820 26936 135620 27056
rect 134820 25848 135620 25968
rect 134820 24896 135620 25016
rect 134820 23808 135620 23928
rect 134820 22856 135620 22976
rect 134820 21768 135620 21888
rect 134820 20816 135620 20936
rect 134820 19728 135620 19848
rect 134820 18776 135620 18896
rect 134820 17688 135620 17808
rect 134820 16736 135620 16856
rect 134820 15648 135620 15768
rect 134820 14696 135620 14816
rect 134820 13608 135620 13728
rect 134820 12656 135620 12776
rect 134820 11568 135620 11688
rect 134820 10616 135620 10736
rect 134820 9528 135620 9648
rect 134820 8576 135620 8696
rect 134820 7488 135620 7608
rect 134820 6536 135620 6656
rect 134820 5448 135620 5568
rect 134820 4496 135620 4616
rect 134820 3408 135620 3528
rect 134820 2456 135620 2576
rect 134820 1368 135620 1488
rect 134820 416 135620 536
<< obsm3 >>
rect 1 133488 134847 134060
rect 1 133208 134740 133488
rect 1 132400 134847 133208
rect 1 132120 134740 132400
rect 1 131448 134847 132120
rect 1 131168 134740 131448
rect 1 130360 134847 131168
rect 1 130080 134740 130360
rect 1 129408 134847 130080
rect 1 129128 134740 129408
rect 1 128320 134847 129128
rect 1 128040 134740 128320
rect 1 127368 134847 128040
rect 1 127088 134740 127368
rect 1 126280 134847 127088
rect 1 126000 134740 126280
rect 1 125328 134847 126000
rect 1 125048 134740 125328
rect 1 124240 134847 125048
rect 1 123960 134740 124240
rect 1 123288 134847 123960
rect 1 123008 134740 123288
rect 1 122200 134847 123008
rect 1 121920 134740 122200
rect 1 121248 134847 121920
rect 1 120968 134740 121248
rect 1 120160 134847 120968
rect 1 119880 134740 120160
rect 1 119208 134847 119880
rect 1 118928 134740 119208
rect 1 118120 134847 118928
rect 1 117840 134740 118120
rect 1 117168 134847 117840
rect 1 116888 134740 117168
rect 1 116080 134847 116888
rect 1 115800 134740 116080
rect 1 115128 134847 115800
rect 1 114848 134740 115128
rect 1 114040 134847 114848
rect 1 113760 134740 114040
rect 1 113088 134847 113760
rect 1 112808 134740 113088
rect 1 112000 134847 112808
rect 1 111720 134740 112000
rect 1 111048 134847 111720
rect 1 110768 134740 111048
rect 1 109960 134847 110768
rect 1 109680 134740 109960
rect 1 108872 134847 109680
rect 1 108592 134740 108872
rect 1 107920 134847 108592
rect 1 107640 134740 107920
rect 1 106832 134847 107640
rect 1 106552 134740 106832
rect 1 105880 134847 106552
rect 1 105600 134740 105880
rect 1 104792 134847 105600
rect 1 104512 134740 104792
rect 1 103840 134847 104512
rect 1 103560 134740 103840
rect 1 102752 134847 103560
rect 1 102472 134740 102752
rect 1 101800 134847 102472
rect 1 101520 134740 101800
rect 1 100712 134847 101520
rect 1 100432 134740 100712
rect 1 99760 134847 100432
rect 1 99480 134740 99760
rect 1 98672 134847 99480
rect 1 98392 134740 98672
rect 1 97720 134847 98392
rect 1 97440 134740 97720
rect 1 96632 134847 97440
rect 1 96352 134740 96632
rect 1 95680 134847 96352
rect 1 95400 134740 95680
rect 1 94592 134847 95400
rect 1 94312 134740 94592
rect 1 93640 134847 94312
rect 1 93360 134740 93640
rect 1 92552 134847 93360
rect 1 92272 134740 92552
rect 1 91600 134847 92272
rect 1 91320 134740 91600
rect 1 90512 134847 91320
rect 1 90232 134740 90512
rect 1 89560 134847 90232
rect 1 89280 134740 89560
rect 1 88472 134847 89280
rect 1 88192 134740 88472
rect 1 87520 134847 88192
rect 1 87240 134740 87520
rect 1 86432 134847 87240
rect 1 86152 134740 86432
rect 1 85480 134847 86152
rect 1 85200 134740 85480
rect 1 84392 134847 85200
rect 1 84112 134740 84392
rect 1 83440 134847 84112
rect 1 83160 134740 83440
rect 1 82352 134847 83160
rect 1 82072 134740 82352
rect 1 81264 134847 82072
rect 1 80984 134740 81264
rect 1 80312 134847 80984
rect 1 80032 134740 80312
rect 1 79224 134847 80032
rect 1 78944 134740 79224
rect 1 78272 134847 78944
rect 1 77992 134740 78272
rect 1 77184 134847 77992
rect 1 76904 134740 77184
rect 1 76232 134847 76904
rect 1 75952 134740 76232
rect 1 75144 134847 75952
rect 1 74864 134740 75144
rect 1 74192 134847 74864
rect 1 73912 134740 74192
rect 1 73104 134847 73912
rect 1 72824 134740 73104
rect 1 72152 134847 72824
rect 1 71872 134740 72152
rect 1 71064 134847 71872
rect 1 70784 134740 71064
rect 1 70112 134847 70784
rect 1 69832 134740 70112
rect 1 69024 134847 69832
rect 1 68744 134740 69024
rect 1 68072 134847 68744
rect 1 67792 134740 68072
rect 1 66984 134847 67792
rect 1 66704 134740 66984
rect 1 66032 134847 66704
rect 1 65752 134740 66032
rect 1 64944 134847 65752
rect 1 64664 134740 64944
rect 1 63992 134847 64664
rect 1 63712 134740 63992
rect 1 62904 134847 63712
rect 1 62624 134740 62904
rect 1 61952 134847 62624
rect 1 61672 134740 61952
rect 1 60864 134847 61672
rect 1 60584 134740 60864
rect 1 59912 134847 60584
rect 1 59632 134740 59912
rect 1 58824 134847 59632
rect 1 58544 134740 58824
rect 1 57872 134847 58544
rect 1 57592 134740 57872
rect 1 56784 134847 57592
rect 1 56504 134740 56784
rect 1 55832 134847 56504
rect 1 55552 134740 55832
rect 1 54744 134847 55552
rect 1 54464 134740 54744
rect 1 53656 134847 54464
rect 1 53376 134740 53656
rect 1 52704 134847 53376
rect 1 52424 134740 52704
rect 1 51616 134847 52424
rect 1 51336 134740 51616
rect 1 50664 134847 51336
rect 1 50384 134740 50664
rect 1 49576 134847 50384
rect 1 49296 134740 49576
rect 1 48624 134847 49296
rect 1 48344 134740 48624
rect 1 47536 134847 48344
rect 1 47256 134740 47536
rect 1 46584 134847 47256
rect 1 46304 134740 46584
rect 1 45496 134847 46304
rect 1 45216 134740 45496
rect 1 44544 134847 45216
rect 1 44264 134740 44544
rect 1 43456 134847 44264
rect 1 43176 134740 43456
rect 1 42504 134847 43176
rect 1 42224 134740 42504
rect 1 41416 134847 42224
rect 1 41136 134740 41416
rect 1 40464 134847 41136
rect 1 40184 134740 40464
rect 1 39376 134847 40184
rect 1 39096 134740 39376
rect 1 38424 134847 39096
rect 1 38144 134740 38424
rect 1 37336 134847 38144
rect 1 37056 134740 37336
rect 1 36384 134847 37056
rect 1 36104 134740 36384
rect 1 35296 134847 36104
rect 1 35016 134740 35296
rect 1 34344 134847 35016
rect 1 34064 134740 34344
rect 1 33256 134847 34064
rect 1 32976 134740 33256
rect 1 32304 134847 32976
rect 1 32024 134740 32304
rect 1 31216 134847 32024
rect 1 30936 134740 31216
rect 1 30264 134847 30936
rect 1 29984 134740 30264
rect 1 29176 134847 29984
rect 1 28896 134740 29176
rect 1 28224 134847 28896
rect 1 27944 134740 28224
rect 1 27136 134847 27944
rect 1 26856 134740 27136
rect 1 26048 134847 26856
rect 1 25768 134740 26048
rect 1 25096 134847 25768
rect 1 24816 134740 25096
rect 1 24008 134847 24816
rect 1 23728 134740 24008
rect 1 23056 134847 23728
rect 1 22776 134740 23056
rect 1 21968 134847 22776
rect 1 21688 134740 21968
rect 1 21016 134847 21688
rect 1 20736 134740 21016
rect 1 19928 134847 20736
rect 1 19648 134740 19928
rect 1 18976 134847 19648
rect 1 18696 134740 18976
rect 1 17888 134847 18696
rect 1 17608 134740 17888
rect 1 16936 134847 17608
rect 1 16656 134740 16936
rect 1 15848 134847 16656
rect 1 15568 134740 15848
rect 1 14896 134847 15568
rect 1 14616 134740 14896
rect 1 13808 134847 14616
rect 1 13528 134740 13808
rect 1 12856 134847 13528
rect 1 12576 134740 12856
rect 1 11768 134847 12576
rect 1 11488 134740 11768
rect 1 10816 134847 11488
rect 1 10536 134740 10816
rect 1 9728 134847 10536
rect 1 9448 134740 9728
rect 1 8776 134847 9448
rect 1 8496 134740 8776
rect 1 7688 134847 8496
rect 1 7408 134740 7688
rect 1 6736 134847 7408
rect 1 6456 134740 6736
rect 1 5648 134847 6456
rect 1 5368 134740 5648
rect 1 4696 134847 5368
rect 1 4416 134740 4696
rect 1 3608 134847 4416
rect 1 3328 134740 3608
rect 1 2656 134847 3328
rect 1 2376 134740 2656
rect 1 1568 134847 2376
rect 1 1288 134740 1568
rect 1 616 134847 1288
rect 1 336 134740 616
rect 1 35 134847 336
<< metal4 >>
rect 3828 2128 4148 133872
rect 4488 2176 4808 133824
rect 5148 2176 5468 133824
rect 5808 2176 6128 133824
rect 19188 2128 19508 133872
rect 19848 2176 20168 133824
rect 20508 2176 20828 133824
rect 21168 2176 21488 133824
rect 34548 2128 34868 133872
rect 35208 2176 35528 133824
rect 35868 2176 36188 133824
rect 36528 2176 36848 133824
rect 49908 2128 50228 133872
rect 50568 2176 50888 133824
rect 51228 2176 51548 133824
rect 51888 2176 52208 133824
rect 65268 2128 65588 133872
rect 65928 2176 66248 133824
rect 66588 2176 66908 133824
rect 67248 2176 67568 133824
rect 80628 2128 80948 133872
rect 81288 2176 81608 133824
rect 81948 2176 82268 133824
rect 82608 2176 82928 133824
rect 95988 2128 96308 133872
rect 96648 2176 96968 133824
rect 97308 2176 97628 133824
rect 97968 2176 98288 133824
rect 111348 2128 111668 133872
rect 112008 2176 112328 133824
rect 112668 2176 112988 133824
rect 113328 2176 113648 133824
rect 126708 2128 127028 133872
rect 127368 2176 127688 133824
rect 128028 2176 128348 133824
rect 128688 2176 129008 133824
<< obsm4 >>
rect 2807 133952 133329 134061
rect 2807 2891 3748 133952
rect 4228 133904 19108 133952
rect 4228 2891 4408 133904
rect 4888 2891 5068 133904
rect 5548 2891 5728 133904
rect 6208 2891 19108 133904
rect 19588 133904 34468 133952
rect 19588 2891 19768 133904
rect 20248 2891 20428 133904
rect 20908 2891 21088 133904
rect 21568 2891 34468 133904
rect 34948 133904 49828 133952
rect 34948 2891 35128 133904
rect 35608 2891 35788 133904
rect 36268 2891 36448 133904
rect 36928 2891 49828 133904
rect 50308 133904 65188 133952
rect 50308 2891 50488 133904
rect 50968 2891 51148 133904
rect 51628 2891 51808 133904
rect 52288 2891 65188 133904
rect 65668 133904 80548 133952
rect 65668 2891 65848 133904
rect 66328 2891 66508 133904
rect 66988 2891 67168 133904
rect 67648 2891 80548 133904
rect 81028 133904 95908 133952
rect 81028 2891 81208 133904
rect 81688 2891 81868 133904
rect 82348 2891 82528 133904
rect 83008 2891 95908 133904
rect 96388 133904 111268 133952
rect 96388 2891 96568 133904
rect 97048 2891 97228 133904
rect 97708 2891 97888 133904
rect 98368 2891 111268 133904
rect 111748 133904 126628 133952
rect 111748 2891 111928 133904
rect 112408 2891 112588 133904
rect 113068 2891 113248 133904
rect 113728 2891 126628 133904
rect 127108 133904 133329 133952
rect 127108 2891 127288 133904
rect 127768 2891 127948 133904
rect 128428 2891 128608 133904
rect 129088 2891 133329 133904
<< labels >>
rlabel metal3 s 134820 416 135620 536 6 clk
port 1 nsew signal input
rlabel metal2 s 132762 0 132818 800 6 flush_in
port 2 nsew signal input
rlabel metal2 s 6 0 62 800 6 i_in[0]
port 3 nsew signal input
rlabel metal2 s 7826 0 7882 800 6 i_in[10]
port 4 nsew signal input
rlabel metal2 s 8562 0 8618 800 6 i_in[11]
port 5 nsew signal input
rlabel metal2 s 9390 0 9446 800 6 i_in[12]
port 6 nsew signal input
rlabel metal2 s 10218 0 10274 800 6 i_in[13]
port 7 nsew signal input
rlabel metal2 s 10954 0 11010 800 6 i_in[14]
port 8 nsew signal input
rlabel metal2 s 11782 0 11838 800 6 i_in[15]
port 9 nsew signal input
rlabel metal2 s 12518 0 12574 800 6 i_in[16]
port 10 nsew signal input
rlabel metal2 s 13346 0 13402 800 6 i_in[17]
port 11 nsew signal input
rlabel metal2 s 14082 0 14138 800 6 i_in[18]
port 12 nsew signal input
rlabel metal2 s 14910 0 14966 800 6 i_in[19]
port 13 nsew signal input
rlabel metal2 s 742 0 798 800 6 i_in[1]
port 14 nsew signal input
rlabel metal2 s 15646 0 15702 800 6 i_in[20]
port 15 nsew signal input
rlabel metal2 s 16474 0 16530 800 6 i_in[21]
port 16 nsew signal input
rlabel metal2 s 17210 0 17266 800 6 i_in[22]
port 17 nsew signal input
rlabel metal2 s 18038 0 18094 800 6 i_in[23]
port 18 nsew signal input
rlabel metal2 s 18866 0 18922 800 6 i_in[24]
port 19 nsew signal input
rlabel metal2 s 19602 0 19658 800 6 i_in[25]
port 20 nsew signal input
rlabel metal2 s 20430 0 20486 800 6 i_in[26]
port 21 nsew signal input
rlabel metal2 s 21166 0 21222 800 6 i_in[27]
port 22 nsew signal input
rlabel metal2 s 21994 0 22050 800 6 i_in[28]
port 23 nsew signal input
rlabel metal2 s 22730 0 22786 800 6 i_in[29]
port 24 nsew signal input
rlabel metal2 s 1570 0 1626 800 6 i_in[2]
port 25 nsew signal input
rlabel metal2 s 23558 0 23614 800 6 i_in[30]
port 26 nsew signal input
rlabel metal2 s 24294 0 24350 800 6 i_in[31]
port 27 nsew signal input
rlabel metal2 s 25122 0 25178 800 6 i_in[32]
port 28 nsew signal input
rlabel metal2 s 25858 0 25914 800 6 i_in[33]
port 29 nsew signal input
rlabel metal2 s 26686 0 26742 800 6 i_in[34]
port 30 nsew signal input
rlabel metal2 s 27514 0 27570 800 6 i_in[35]
port 31 nsew signal input
rlabel metal2 s 28250 0 28306 800 6 i_in[36]
port 32 nsew signal input
rlabel metal2 s 29078 0 29134 800 6 i_in[37]
port 33 nsew signal input
rlabel metal2 s 29814 0 29870 800 6 i_in[38]
port 34 nsew signal input
rlabel metal2 s 30642 0 30698 800 6 i_in[39]
port 35 nsew signal input
rlabel metal2 s 2306 0 2362 800 6 i_in[3]
port 36 nsew signal input
rlabel metal2 s 31378 0 31434 800 6 i_in[40]
port 37 nsew signal input
rlabel metal2 s 32206 0 32262 800 6 i_in[41]
port 38 nsew signal input
rlabel metal2 s 32942 0 32998 800 6 i_in[42]
port 39 nsew signal input
rlabel metal2 s 33770 0 33826 800 6 i_in[43]
port 40 nsew signal input
rlabel metal2 s 34506 0 34562 800 6 i_in[44]
port 41 nsew signal input
rlabel metal2 s 35334 0 35390 800 6 i_in[45]
port 42 nsew signal input
rlabel metal2 s 36070 0 36126 800 6 i_in[46]
port 43 nsew signal input
rlabel metal2 s 36898 0 36954 800 6 i_in[47]
port 44 nsew signal input
rlabel metal2 s 37726 0 37782 800 6 i_in[48]
port 45 nsew signal input
rlabel metal2 s 38462 0 38518 800 6 i_in[49]
port 46 nsew signal input
rlabel metal2 s 3134 0 3190 800 6 i_in[4]
port 47 nsew signal input
rlabel metal2 s 39290 0 39346 800 6 i_in[50]
port 48 nsew signal input
rlabel metal2 s 40026 0 40082 800 6 i_in[51]
port 49 nsew signal input
rlabel metal2 s 40854 0 40910 800 6 i_in[52]
port 50 nsew signal input
rlabel metal2 s 41590 0 41646 800 6 i_in[53]
port 51 nsew signal input
rlabel metal2 s 42418 0 42474 800 6 i_in[54]
port 52 nsew signal input
rlabel metal2 s 43154 0 43210 800 6 i_in[55]
port 53 nsew signal input
rlabel metal2 s 43982 0 44038 800 6 i_in[56]
port 54 nsew signal input
rlabel metal2 s 44718 0 44774 800 6 i_in[57]
port 55 nsew signal input
rlabel metal2 s 45546 0 45602 800 6 i_in[58]
port 56 nsew signal input
rlabel metal2 s 46374 0 46430 800 6 i_in[59]
port 57 nsew signal input
rlabel metal2 s 3870 0 3926 800 6 i_in[5]
port 58 nsew signal input
rlabel metal2 s 47110 0 47166 800 6 i_in[60]
port 59 nsew signal input
rlabel metal2 s 47938 0 47994 800 6 i_in[61]
port 60 nsew signal input
rlabel metal2 s 48674 0 48730 800 6 i_in[62]
port 61 nsew signal input
rlabel metal2 s 49502 0 49558 800 6 i_in[63]
port 62 nsew signal input
rlabel metal2 s 50238 0 50294 800 6 i_in[64]
port 63 nsew signal input
rlabel metal2 s 51066 0 51122 800 6 i_in[65]
port 64 nsew signal input
rlabel metal2 s 51802 0 51858 800 6 i_in[66]
port 65 nsew signal input
rlabel metal2 s 52630 0 52686 800 6 i_in[67]
port 66 nsew signal input
rlabel metal2 s 53366 0 53422 800 6 i_in[68]
port 67 nsew signal input
rlabel metal2 s 54194 0 54250 800 6 i_in[69]
port 68 nsew signal input
rlabel metal2 s 4698 0 4754 800 6 i_in[6]
port 69 nsew signal input
rlabel metal2 s 5434 0 5490 800 6 i_in[7]
port 70 nsew signal input
rlabel metal2 s 6262 0 6318 800 6 i_in[8]
port 71 nsew signal input
rlabel metal2 s 6998 0 7054 800 6 i_in[9]
port 72 nsew signal input
rlabel metal2 s 55022 0 55078 800 6 i_out[0]
port 73 nsew signal output
rlabel metal2 s 62842 0 62898 800 6 i_out[10]
port 74 nsew signal output
rlabel metal2 s 63670 0 63726 800 6 i_out[11]
port 75 nsew signal output
rlabel metal2 s 64406 0 64462 800 6 i_out[12]
port 76 nsew signal output
rlabel metal2 s 65234 0 65290 800 6 i_out[13]
port 77 nsew signal output
rlabel metal2 s 65970 0 66026 800 6 i_out[14]
port 78 nsew signal output
rlabel metal2 s 66798 0 66854 800 6 i_out[15]
port 79 nsew signal output
rlabel metal2 s 67534 0 67590 800 6 i_out[16]
port 80 nsew signal output
rlabel metal2 s 68362 0 68418 800 6 i_out[17]
port 81 nsew signal output
rlabel metal2 s 69098 0 69154 800 6 i_out[18]
port 82 nsew signal output
rlabel metal2 s 69926 0 69982 800 6 i_out[19]
port 83 nsew signal output
rlabel metal2 s 55758 0 55814 800 6 i_out[1]
port 84 nsew signal output
rlabel metal2 s 70662 0 70718 800 6 i_out[20]
port 85 nsew signal output
rlabel metal2 s 71490 0 71546 800 6 i_out[21]
port 86 nsew signal output
rlabel metal2 s 72226 0 72282 800 6 i_out[22]
port 87 nsew signal output
rlabel metal2 s 73054 0 73110 800 6 i_out[23]
port 88 nsew signal output
rlabel metal2 s 73882 0 73938 800 6 i_out[24]
port 89 nsew signal output
rlabel metal2 s 74618 0 74674 800 6 i_out[25]
port 90 nsew signal output
rlabel metal2 s 75446 0 75502 800 6 i_out[26]
port 91 nsew signal output
rlabel metal2 s 76182 0 76238 800 6 i_out[27]
port 92 nsew signal output
rlabel metal2 s 77010 0 77066 800 6 i_out[28]
port 93 nsew signal output
rlabel metal2 s 77746 0 77802 800 6 i_out[29]
port 94 nsew signal output
rlabel metal2 s 56586 0 56642 800 6 i_out[2]
port 95 nsew signal output
rlabel metal2 s 78574 0 78630 800 6 i_out[30]
port 96 nsew signal output
rlabel metal2 s 79310 0 79366 800 6 i_out[31]
port 97 nsew signal output
rlabel metal2 s 80138 0 80194 800 6 i_out[32]
port 98 nsew signal output
rlabel metal2 s 80874 0 80930 800 6 i_out[33]
port 99 nsew signal output
rlabel metal2 s 81702 0 81758 800 6 i_out[34]
port 100 nsew signal output
rlabel metal2 s 82530 0 82586 800 6 i_out[35]
port 101 nsew signal output
rlabel metal2 s 83266 0 83322 800 6 i_out[36]
port 102 nsew signal output
rlabel metal2 s 84094 0 84150 800 6 i_out[37]
port 103 nsew signal output
rlabel metal2 s 84830 0 84886 800 6 i_out[38]
port 104 nsew signal output
rlabel metal2 s 85658 0 85714 800 6 i_out[39]
port 105 nsew signal output
rlabel metal2 s 57322 0 57378 800 6 i_out[3]
port 106 nsew signal output
rlabel metal2 s 86394 0 86450 800 6 i_out[40]
port 107 nsew signal output
rlabel metal2 s 87222 0 87278 800 6 i_out[41]
port 108 nsew signal output
rlabel metal2 s 87958 0 88014 800 6 i_out[42]
port 109 nsew signal output
rlabel metal2 s 88786 0 88842 800 6 i_out[43]
port 110 nsew signal output
rlabel metal2 s 89522 0 89578 800 6 i_out[44]
port 111 nsew signal output
rlabel metal2 s 90350 0 90406 800 6 i_out[45]
port 112 nsew signal output
rlabel metal2 s 91178 0 91234 800 6 i_out[46]
port 113 nsew signal output
rlabel metal2 s 91914 0 91970 800 6 i_out[47]
port 114 nsew signal output
rlabel metal2 s 92742 0 92798 800 6 i_out[48]
port 115 nsew signal output
rlabel metal2 s 93478 0 93534 800 6 i_out[49]
port 116 nsew signal output
rlabel metal2 s 58150 0 58206 800 6 i_out[4]
port 117 nsew signal output
rlabel metal2 s 94306 0 94362 800 6 i_out[50]
port 118 nsew signal output
rlabel metal2 s 95042 0 95098 800 6 i_out[51]
port 119 nsew signal output
rlabel metal2 s 95870 0 95926 800 6 i_out[52]
port 120 nsew signal output
rlabel metal2 s 96606 0 96662 800 6 i_out[53]
port 121 nsew signal output
rlabel metal2 s 97434 0 97490 800 6 i_out[54]
port 122 nsew signal output
rlabel metal2 s 98170 0 98226 800 6 i_out[55]
port 123 nsew signal output
rlabel metal2 s 98998 0 99054 800 6 i_out[56]
port 124 nsew signal output
rlabel metal2 s 99826 0 99882 800 6 i_out[57]
port 125 nsew signal output
rlabel metal2 s 100562 0 100618 800 6 i_out[58]
port 126 nsew signal output
rlabel metal2 s 101390 0 101446 800 6 i_out[59]
port 127 nsew signal output
rlabel metal2 s 58886 0 58942 800 6 i_out[5]
port 128 nsew signal output
rlabel metal2 s 102126 0 102182 800 6 i_out[60]
port 129 nsew signal output
rlabel metal2 s 102954 0 103010 800 6 i_out[61]
port 130 nsew signal output
rlabel metal2 s 103690 0 103746 800 6 i_out[62]
port 131 nsew signal output
rlabel metal2 s 104518 0 104574 800 6 i_out[63]
port 132 nsew signal output
rlabel metal2 s 105254 0 105310 800 6 i_out[64]
port 133 nsew signal output
rlabel metal2 s 106082 0 106138 800 6 i_out[65]
port 134 nsew signal output
rlabel metal2 s 106818 0 106874 800 6 i_out[66]
port 135 nsew signal output
rlabel metal2 s 107646 0 107702 800 6 i_out[67]
port 136 nsew signal output
rlabel metal2 s 108382 0 108438 800 6 i_out[68]
port 137 nsew signal output
rlabel metal2 s 109210 0 109266 800 6 i_out[69]
port 138 nsew signal output
rlabel metal2 s 59714 0 59770 800 6 i_out[6]
port 139 nsew signal output
rlabel metal2 s 110038 0 110094 800 6 i_out[70]
port 140 nsew signal output
rlabel metal2 s 110774 0 110830 800 6 i_out[71]
port 141 nsew signal output
rlabel metal2 s 111602 0 111658 800 6 i_out[72]
port 142 nsew signal output
rlabel metal2 s 112338 0 112394 800 6 i_out[73]
port 143 nsew signal output
rlabel metal2 s 113166 0 113222 800 6 i_out[74]
port 144 nsew signal output
rlabel metal2 s 113902 0 113958 800 6 i_out[75]
port 145 nsew signal output
rlabel metal2 s 114730 0 114786 800 6 i_out[76]
port 146 nsew signal output
rlabel metal2 s 115466 0 115522 800 6 i_out[77]
port 147 nsew signal output
rlabel metal2 s 116294 0 116350 800 6 i_out[78]
port 148 nsew signal output
rlabel metal2 s 117030 0 117086 800 6 i_out[79]
port 149 nsew signal output
rlabel metal2 s 60450 0 60506 800 6 i_out[7]
port 150 nsew signal output
rlabel metal2 s 117858 0 117914 800 6 i_out[80]
port 151 nsew signal output
rlabel metal2 s 118686 0 118742 800 6 i_out[81]
port 152 nsew signal output
rlabel metal2 s 119422 0 119478 800 6 i_out[82]
port 153 nsew signal output
rlabel metal2 s 120250 0 120306 800 6 i_out[83]
port 154 nsew signal output
rlabel metal2 s 120986 0 121042 800 6 i_out[84]
port 155 nsew signal output
rlabel metal2 s 121814 0 121870 800 6 i_out[85]
port 156 nsew signal output
rlabel metal2 s 122550 0 122606 800 6 i_out[86]
port 157 nsew signal output
rlabel metal2 s 123378 0 123434 800 6 i_out[87]
port 158 nsew signal output
rlabel metal2 s 124114 0 124170 800 6 i_out[88]
port 159 nsew signal output
rlabel metal2 s 124942 0 124998 800 6 i_out[89]
port 160 nsew signal output
rlabel metal2 s 61278 0 61334 800 6 i_out[8]
port 161 nsew signal output
rlabel metal2 s 125678 0 125734 800 6 i_out[90]
port 162 nsew signal output
rlabel metal2 s 126506 0 126562 800 6 i_out[91]
port 163 nsew signal output
rlabel metal2 s 127334 0 127390 800 6 i_out[92]
port 164 nsew signal output
rlabel metal2 s 128070 0 128126 800 6 i_out[93]
port 165 nsew signal output
rlabel metal2 s 128898 0 128954 800 6 i_out[94]
port 166 nsew signal output
rlabel metal2 s 129634 0 129690 800 6 i_out[95]
port 167 nsew signal output
rlabel metal2 s 130462 0 130518 800 6 i_out[96]
port 168 nsew signal output
rlabel metal2 s 131198 0 131254 800 6 i_out[97]
port 169 nsew signal output
rlabel metal2 s 132026 0 132082 800 6 i_out[98]
port 170 nsew signal output
rlabel metal2 s 62014 0 62070 800 6 i_out[9]
port 171 nsew signal output
rlabel metal2 s 133590 0 133646 800 6 inval_in
port 172 nsew signal input
rlabel metal3 s 134820 2456 135620 2576 6 m_in[0]
port 173 nsew signal input
rlabel metal3 s 134820 104592 135620 104712 6 m_in[100]
port 174 nsew signal input
rlabel metal3 s 134820 105680 135620 105800 6 m_in[101]
port 175 nsew signal input
rlabel metal3 s 134820 106632 135620 106752 6 m_in[102]
port 176 nsew signal input
rlabel metal3 s 134820 107720 135620 107840 6 m_in[103]
port 177 nsew signal input
rlabel metal3 s 134820 108672 135620 108792 6 m_in[104]
port 178 nsew signal input
rlabel metal3 s 134820 109760 135620 109880 6 m_in[105]
port 179 nsew signal input
rlabel metal3 s 134820 110848 135620 110968 6 m_in[106]
port 180 nsew signal input
rlabel metal3 s 134820 111800 135620 111920 6 m_in[107]
port 181 nsew signal input
rlabel metal3 s 134820 112888 135620 113008 6 m_in[108]
port 182 nsew signal input
rlabel metal3 s 134820 113840 135620 113960 6 m_in[109]
port 183 nsew signal input
rlabel metal3 s 134820 12656 135620 12776 6 m_in[10]
port 184 nsew signal input
rlabel metal3 s 134820 114928 135620 115048 6 m_in[110]
port 185 nsew signal input
rlabel metal3 s 134820 115880 135620 116000 6 m_in[111]
port 186 nsew signal input
rlabel metal3 s 134820 116968 135620 117088 6 m_in[112]
port 187 nsew signal input
rlabel metal3 s 134820 117920 135620 118040 6 m_in[113]
port 188 nsew signal input
rlabel metal3 s 134820 119008 135620 119128 6 m_in[114]
port 189 nsew signal input
rlabel metal3 s 134820 119960 135620 120080 6 m_in[115]
port 190 nsew signal input
rlabel metal3 s 134820 121048 135620 121168 6 m_in[116]
port 191 nsew signal input
rlabel metal3 s 134820 122000 135620 122120 6 m_in[117]
port 192 nsew signal input
rlabel metal3 s 134820 123088 135620 123208 6 m_in[118]
port 193 nsew signal input
rlabel metal3 s 134820 124040 135620 124160 6 m_in[119]
port 194 nsew signal input
rlabel metal3 s 134820 13608 135620 13728 6 m_in[11]
port 195 nsew signal input
rlabel metal3 s 134820 125128 135620 125248 6 m_in[120]
port 196 nsew signal input
rlabel metal3 s 134820 126080 135620 126200 6 m_in[121]
port 197 nsew signal input
rlabel metal3 s 134820 127168 135620 127288 6 m_in[122]
port 198 nsew signal input
rlabel metal3 s 134820 128120 135620 128240 6 m_in[123]
port 199 nsew signal input
rlabel metal3 s 134820 129208 135620 129328 6 m_in[124]
port 200 nsew signal input
rlabel metal3 s 134820 130160 135620 130280 6 m_in[125]
port 201 nsew signal input
rlabel metal3 s 134820 131248 135620 131368 6 m_in[126]
port 202 nsew signal input
rlabel metal3 s 134820 132200 135620 132320 6 m_in[127]
port 203 nsew signal input
rlabel metal3 s 134820 133288 135620 133408 6 m_in[128]
port 204 nsew signal input
rlabel metal3 s 134820 134240 135620 134360 6 m_in[129]
port 205 nsew signal input
rlabel metal3 s 134820 14696 135620 14816 6 m_in[12]
port 206 nsew signal input
rlabel metal3 s 134820 135328 135620 135448 6 m_in[130]
port 207 nsew signal input
rlabel metal3 s 134820 15648 135620 15768 6 m_in[13]
port 208 nsew signal input
rlabel metal3 s 134820 16736 135620 16856 6 m_in[14]
port 209 nsew signal input
rlabel metal3 s 134820 17688 135620 17808 6 m_in[15]
port 210 nsew signal input
rlabel metal3 s 134820 18776 135620 18896 6 m_in[16]
port 211 nsew signal input
rlabel metal3 s 134820 19728 135620 19848 6 m_in[17]
port 212 nsew signal input
rlabel metal3 s 134820 20816 135620 20936 6 m_in[18]
port 213 nsew signal input
rlabel metal3 s 134820 21768 135620 21888 6 m_in[19]
port 214 nsew signal input
rlabel metal3 s 134820 3408 135620 3528 6 m_in[1]
port 215 nsew signal input
rlabel metal3 s 134820 22856 135620 22976 6 m_in[20]
port 216 nsew signal input
rlabel metal3 s 134820 23808 135620 23928 6 m_in[21]
port 217 nsew signal input
rlabel metal3 s 134820 24896 135620 25016 6 m_in[22]
port 218 nsew signal input
rlabel metal3 s 134820 25848 135620 25968 6 m_in[23]
port 219 nsew signal input
rlabel metal3 s 134820 26936 135620 27056 6 m_in[24]
port 220 nsew signal input
rlabel metal3 s 134820 28024 135620 28144 6 m_in[25]
port 221 nsew signal input
rlabel metal3 s 134820 28976 135620 29096 6 m_in[26]
port 222 nsew signal input
rlabel metal3 s 134820 30064 135620 30184 6 m_in[27]
port 223 nsew signal input
rlabel metal3 s 134820 31016 135620 31136 6 m_in[28]
port 224 nsew signal input
rlabel metal3 s 134820 32104 135620 32224 6 m_in[29]
port 225 nsew signal input
rlabel metal3 s 134820 4496 135620 4616 6 m_in[2]
port 226 nsew signal input
rlabel metal3 s 134820 33056 135620 33176 6 m_in[30]
port 227 nsew signal input
rlabel metal3 s 134820 34144 135620 34264 6 m_in[31]
port 228 nsew signal input
rlabel metal3 s 134820 35096 135620 35216 6 m_in[32]
port 229 nsew signal input
rlabel metal3 s 134820 36184 135620 36304 6 m_in[33]
port 230 nsew signal input
rlabel metal3 s 134820 37136 135620 37256 6 m_in[34]
port 231 nsew signal input
rlabel metal3 s 134820 38224 135620 38344 6 m_in[35]
port 232 nsew signal input
rlabel metal3 s 134820 39176 135620 39296 6 m_in[36]
port 233 nsew signal input
rlabel metal3 s 134820 40264 135620 40384 6 m_in[37]
port 234 nsew signal input
rlabel metal3 s 134820 41216 135620 41336 6 m_in[38]
port 235 nsew signal input
rlabel metal3 s 134820 42304 135620 42424 6 m_in[39]
port 236 nsew signal input
rlabel metal3 s 134820 5448 135620 5568 6 m_in[3]
port 237 nsew signal input
rlabel metal3 s 134820 43256 135620 43376 6 m_in[40]
port 238 nsew signal input
rlabel metal3 s 134820 44344 135620 44464 6 m_in[41]
port 239 nsew signal input
rlabel metal3 s 134820 45296 135620 45416 6 m_in[42]
port 240 nsew signal input
rlabel metal3 s 134820 46384 135620 46504 6 m_in[43]
port 241 nsew signal input
rlabel metal3 s 134820 47336 135620 47456 6 m_in[44]
port 242 nsew signal input
rlabel metal3 s 134820 48424 135620 48544 6 m_in[45]
port 243 nsew signal input
rlabel metal3 s 134820 49376 135620 49496 6 m_in[46]
port 244 nsew signal input
rlabel metal3 s 134820 50464 135620 50584 6 m_in[47]
port 245 nsew signal input
rlabel metal3 s 134820 51416 135620 51536 6 m_in[48]
port 246 nsew signal input
rlabel metal3 s 134820 52504 135620 52624 6 m_in[49]
port 247 nsew signal input
rlabel metal3 s 134820 6536 135620 6656 6 m_in[4]
port 248 nsew signal input
rlabel metal3 s 134820 53456 135620 53576 6 m_in[50]
port 249 nsew signal input
rlabel metal3 s 134820 54544 135620 54664 6 m_in[51]
port 250 nsew signal input
rlabel metal3 s 134820 55632 135620 55752 6 m_in[52]
port 251 nsew signal input
rlabel metal3 s 134820 56584 135620 56704 6 m_in[53]
port 252 nsew signal input
rlabel metal3 s 134820 57672 135620 57792 6 m_in[54]
port 253 nsew signal input
rlabel metal3 s 134820 58624 135620 58744 6 m_in[55]
port 254 nsew signal input
rlabel metal3 s 134820 59712 135620 59832 6 m_in[56]
port 255 nsew signal input
rlabel metal3 s 134820 60664 135620 60784 6 m_in[57]
port 256 nsew signal input
rlabel metal3 s 134820 61752 135620 61872 6 m_in[58]
port 257 nsew signal input
rlabel metal3 s 134820 62704 135620 62824 6 m_in[59]
port 258 nsew signal input
rlabel metal3 s 134820 7488 135620 7608 6 m_in[5]
port 259 nsew signal input
rlabel metal3 s 134820 63792 135620 63912 6 m_in[60]
port 260 nsew signal input
rlabel metal3 s 134820 64744 135620 64864 6 m_in[61]
port 261 nsew signal input
rlabel metal3 s 134820 65832 135620 65952 6 m_in[62]
port 262 nsew signal input
rlabel metal3 s 134820 66784 135620 66904 6 m_in[63]
port 263 nsew signal input
rlabel metal3 s 134820 67872 135620 67992 6 m_in[64]
port 264 nsew signal input
rlabel metal3 s 134820 68824 135620 68944 6 m_in[65]
port 265 nsew signal input
rlabel metal3 s 134820 69912 135620 70032 6 m_in[66]
port 266 nsew signal input
rlabel metal3 s 134820 70864 135620 70984 6 m_in[67]
port 267 nsew signal input
rlabel metal3 s 134820 71952 135620 72072 6 m_in[68]
port 268 nsew signal input
rlabel metal3 s 134820 72904 135620 73024 6 m_in[69]
port 269 nsew signal input
rlabel metal3 s 134820 8576 135620 8696 6 m_in[6]
port 270 nsew signal input
rlabel metal3 s 134820 73992 135620 74112 6 m_in[70]
port 271 nsew signal input
rlabel metal3 s 134820 74944 135620 75064 6 m_in[71]
port 272 nsew signal input
rlabel metal3 s 134820 76032 135620 76152 6 m_in[72]
port 273 nsew signal input
rlabel metal3 s 134820 76984 135620 77104 6 m_in[73]
port 274 nsew signal input
rlabel metal3 s 134820 78072 135620 78192 6 m_in[74]
port 275 nsew signal input
rlabel metal3 s 134820 79024 135620 79144 6 m_in[75]
port 276 nsew signal input
rlabel metal3 s 134820 80112 135620 80232 6 m_in[76]
port 277 nsew signal input
rlabel metal3 s 134820 81064 135620 81184 6 m_in[77]
port 278 nsew signal input
rlabel metal3 s 134820 82152 135620 82272 6 m_in[78]
port 279 nsew signal input
rlabel metal3 s 134820 83240 135620 83360 6 m_in[79]
port 280 nsew signal input
rlabel metal3 s 134820 9528 135620 9648 6 m_in[7]
port 281 nsew signal input
rlabel metal3 s 134820 84192 135620 84312 6 m_in[80]
port 282 nsew signal input
rlabel metal3 s 134820 85280 135620 85400 6 m_in[81]
port 283 nsew signal input
rlabel metal3 s 134820 86232 135620 86352 6 m_in[82]
port 284 nsew signal input
rlabel metal3 s 134820 87320 135620 87440 6 m_in[83]
port 285 nsew signal input
rlabel metal3 s 134820 88272 135620 88392 6 m_in[84]
port 286 nsew signal input
rlabel metal3 s 134820 89360 135620 89480 6 m_in[85]
port 287 nsew signal input
rlabel metal3 s 134820 90312 135620 90432 6 m_in[86]
port 288 nsew signal input
rlabel metal3 s 134820 91400 135620 91520 6 m_in[87]
port 289 nsew signal input
rlabel metal3 s 134820 92352 135620 92472 6 m_in[88]
port 290 nsew signal input
rlabel metal3 s 134820 93440 135620 93560 6 m_in[89]
port 291 nsew signal input
rlabel metal3 s 134820 10616 135620 10736 6 m_in[8]
port 292 nsew signal input
rlabel metal3 s 134820 94392 135620 94512 6 m_in[90]
port 293 nsew signal input
rlabel metal3 s 134820 95480 135620 95600 6 m_in[91]
port 294 nsew signal input
rlabel metal3 s 134820 96432 135620 96552 6 m_in[92]
port 295 nsew signal input
rlabel metal3 s 134820 97520 135620 97640 6 m_in[93]
port 296 nsew signal input
rlabel metal3 s 134820 98472 135620 98592 6 m_in[94]
port 297 nsew signal input
rlabel metal3 s 134820 99560 135620 99680 6 m_in[95]
port 298 nsew signal input
rlabel metal3 s 134820 100512 135620 100632 6 m_in[96]
port 299 nsew signal input
rlabel metal3 s 134820 101600 135620 101720 6 m_in[97]
port 300 nsew signal input
rlabel metal3 s 134820 102552 135620 102672 6 m_in[98]
port 301 nsew signal input
rlabel metal3 s 134820 103640 135620 103760 6 m_in[99]
port 302 nsew signal input
rlabel metal3 s 134820 11568 135620 11688 6 m_in[9]
port 303 nsew signal input
rlabel metal3 s 134820 1368 135620 1488 6 rst
port 304 nsew signal input
rlabel metal2 s 134326 0 134382 800 6 stall_in
port 305 nsew signal input
rlabel metal2 s 135154 0 135210 800 6 stall_out
port 306 nsew signal output
rlabel metal2 s 6 135200 62 136000 6 wishbone_in[0]
port 307 nsew signal input
rlabel metal2 s 7826 135200 7882 136000 6 wishbone_in[10]
port 308 nsew signal input
rlabel metal2 s 8562 135200 8618 136000 6 wishbone_in[11]
port 309 nsew signal input
rlabel metal2 s 9390 135200 9446 136000 6 wishbone_in[12]
port 310 nsew signal input
rlabel metal2 s 10218 135200 10274 136000 6 wishbone_in[13]
port 311 nsew signal input
rlabel metal2 s 10954 135200 11010 136000 6 wishbone_in[14]
port 312 nsew signal input
rlabel metal2 s 11782 135200 11838 136000 6 wishbone_in[15]
port 313 nsew signal input
rlabel metal2 s 12518 135200 12574 136000 6 wishbone_in[16]
port 314 nsew signal input
rlabel metal2 s 13346 135200 13402 136000 6 wishbone_in[17]
port 315 nsew signal input
rlabel metal2 s 14082 135200 14138 136000 6 wishbone_in[18]
port 316 nsew signal input
rlabel metal2 s 14910 135200 14966 136000 6 wishbone_in[19]
port 317 nsew signal input
rlabel metal2 s 742 135200 798 136000 6 wishbone_in[1]
port 318 nsew signal input
rlabel metal2 s 15646 135200 15702 136000 6 wishbone_in[20]
port 319 nsew signal input
rlabel metal2 s 16474 135200 16530 136000 6 wishbone_in[21]
port 320 nsew signal input
rlabel metal2 s 17210 135200 17266 136000 6 wishbone_in[22]
port 321 nsew signal input
rlabel metal2 s 18038 135200 18094 136000 6 wishbone_in[23]
port 322 nsew signal input
rlabel metal2 s 18866 135200 18922 136000 6 wishbone_in[24]
port 323 nsew signal input
rlabel metal2 s 19602 135200 19658 136000 6 wishbone_in[25]
port 324 nsew signal input
rlabel metal2 s 20430 135200 20486 136000 6 wishbone_in[26]
port 325 nsew signal input
rlabel metal2 s 21166 135200 21222 136000 6 wishbone_in[27]
port 326 nsew signal input
rlabel metal2 s 21994 135200 22050 136000 6 wishbone_in[28]
port 327 nsew signal input
rlabel metal2 s 22730 135200 22786 136000 6 wishbone_in[29]
port 328 nsew signal input
rlabel metal2 s 1570 135200 1626 136000 6 wishbone_in[2]
port 329 nsew signal input
rlabel metal2 s 23558 135200 23614 136000 6 wishbone_in[30]
port 330 nsew signal input
rlabel metal2 s 24294 135200 24350 136000 6 wishbone_in[31]
port 331 nsew signal input
rlabel metal2 s 25122 135200 25178 136000 6 wishbone_in[32]
port 332 nsew signal input
rlabel metal2 s 25858 135200 25914 136000 6 wishbone_in[33]
port 333 nsew signal input
rlabel metal2 s 26686 135200 26742 136000 6 wishbone_in[34]
port 334 nsew signal input
rlabel metal2 s 27514 135200 27570 136000 6 wishbone_in[35]
port 335 nsew signal input
rlabel metal2 s 28250 135200 28306 136000 6 wishbone_in[36]
port 336 nsew signal input
rlabel metal2 s 29078 135200 29134 136000 6 wishbone_in[37]
port 337 nsew signal input
rlabel metal2 s 29814 135200 29870 136000 6 wishbone_in[38]
port 338 nsew signal input
rlabel metal2 s 30642 135200 30698 136000 6 wishbone_in[39]
port 339 nsew signal input
rlabel metal2 s 2306 135200 2362 136000 6 wishbone_in[3]
port 340 nsew signal input
rlabel metal2 s 31378 135200 31434 136000 6 wishbone_in[40]
port 341 nsew signal input
rlabel metal2 s 32206 135200 32262 136000 6 wishbone_in[41]
port 342 nsew signal input
rlabel metal2 s 32942 135200 32998 136000 6 wishbone_in[42]
port 343 nsew signal input
rlabel metal2 s 33770 135200 33826 136000 6 wishbone_in[43]
port 344 nsew signal input
rlabel metal2 s 34506 135200 34562 136000 6 wishbone_in[44]
port 345 nsew signal input
rlabel metal2 s 35334 135200 35390 136000 6 wishbone_in[45]
port 346 nsew signal input
rlabel metal2 s 36070 135200 36126 136000 6 wishbone_in[46]
port 347 nsew signal input
rlabel metal2 s 36898 135200 36954 136000 6 wishbone_in[47]
port 348 nsew signal input
rlabel metal2 s 37726 135200 37782 136000 6 wishbone_in[48]
port 349 nsew signal input
rlabel metal2 s 38462 135200 38518 136000 6 wishbone_in[49]
port 350 nsew signal input
rlabel metal2 s 3134 135200 3190 136000 6 wishbone_in[4]
port 351 nsew signal input
rlabel metal2 s 39290 135200 39346 136000 6 wishbone_in[50]
port 352 nsew signal input
rlabel metal2 s 40026 135200 40082 136000 6 wishbone_in[51]
port 353 nsew signal input
rlabel metal2 s 40854 135200 40910 136000 6 wishbone_in[52]
port 354 nsew signal input
rlabel metal2 s 41590 135200 41646 136000 6 wishbone_in[53]
port 355 nsew signal input
rlabel metal2 s 42418 135200 42474 136000 6 wishbone_in[54]
port 356 nsew signal input
rlabel metal2 s 43154 135200 43210 136000 6 wishbone_in[55]
port 357 nsew signal input
rlabel metal2 s 43982 135200 44038 136000 6 wishbone_in[56]
port 358 nsew signal input
rlabel metal2 s 44718 135200 44774 136000 6 wishbone_in[57]
port 359 nsew signal input
rlabel metal2 s 45546 135200 45602 136000 6 wishbone_in[58]
port 360 nsew signal input
rlabel metal2 s 46374 135200 46430 136000 6 wishbone_in[59]
port 361 nsew signal input
rlabel metal2 s 3870 135200 3926 136000 6 wishbone_in[5]
port 362 nsew signal input
rlabel metal2 s 47110 135200 47166 136000 6 wishbone_in[60]
port 363 nsew signal input
rlabel metal2 s 47938 135200 47994 136000 6 wishbone_in[61]
port 364 nsew signal input
rlabel metal2 s 48674 135200 48730 136000 6 wishbone_in[62]
port 365 nsew signal input
rlabel metal2 s 49502 135200 49558 136000 6 wishbone_in[63]
port 366 nsew signal input
rlabel metal2 s 50238 135200 50294 136000 6 wishbone_in[64]
port 367 nsew signal input
rlabel metal2 s 51066 135200 51122 136000 6 wishbone_in[65]
port 368 nsew signal input
rlabel metal2 s 4698 135200 4754 136000 6 wishbone_in[6]
port 369 nsew signal input
rlabel metal2 s 5434 135200 5490 136000 6 wishbone_in[7]
port 370 nsew signal input
rlabel metal2 s 6262 135200 6318 136000 6 wishbone_in[8]
port 371 nsew signal input
rlabel metal2 s 6998 135200 7054 136000 6 wishbone_in[9]
port 372 nsew signal input
rlabel metal2 s 51802 135200 51858 136000 6 wishbone_out[0]
port 373 nsew signal output
rlabel metal2 s 130462 135200 130518 136000 6 wishbone_out[100]
port 374 nsew signal output
rlabel metal2 s 131198 135200 131254 136000 6 wishbone_out[101]
port 375 nsew signal output
rlabel metal2 s 132026 135200 132082 136000 6 wishbone_out[102]
port 376 nsew signal output
rlabel metal2 s 132762 135200 132818 136000 6 wishbone_out[103]
port 377 nsew signal output
rlabel metal2 s 133590 135200 133646 136000 6 wishbone_out[104]
port 378 nsew signal output
rlabel metal2 s 134326 135200 134382 136000 6 wishbone_out[105]
port 379 nsew signal output
rlabel metal2 s 135154 135200 135210 136000 6 wishbone_out[106]
port 380 nsew signal output
rlabel metal2 s 59714 135200 59770 136000 6 wishbone_out[10]
port 381 nsew signal output
rlabel metal2 s 60450 135200 60506 136000 6 wishbone_out[11]
port 382 nsew signal output
rlabel metal2 s 61278 135200 61334 136000 6 wishbone_out[12]
port 383 nsew signal output
rlabel metal2 s 62014 135200 62070 136000 6 wishbone_out[13]
port 384 nsew signal output
rlabel metal2 s 62842 135200 62898 136000 6 wishbone_out[14]
port 385 nsew signal output
rlabel metal2 s 63670 135200 63726 136000 6 wishbone_out[15]
port 386 nsew signal output
rlabel metal2 s 64406 135200 64462 136000 6 wishbone_out[16]
port 387 nsew signal output
rlabel metal2 s 65234 135200 65290 136000 6 wishbone_out[17]
port 388 nsew signal output
rlabel metal2 s 65970 135200 66026 136000 6 wishbone_out[18]
port 389 nsew signal output
rlabel metal2 s 66798 135200 66854 136000 6 wishbone_out[19]
port 390 nsew signal output
rlabel metal2 s 52630 135200 52686 136000 6 wishbone_out[1]
port 391 nsew signal output
rlabel metal2 s 67534 135200 67590 136000 6 wishbone_out[20]
port 392 nsew signal output
rlabel metal2 s 68362 135200 68418 136000 6 wishbone_out[21]
port 393 nsew signal output
rlabel metal2 s 69098 135200 69154 136000 6 wishbone_out[22]
port 394 nsew signal output
rlabel metal2 s 69926 135200 69982 136000 6 wishbone_out[23]
port 395 nsew signal output
rlabel metal2 s 70662 135200 70718 136000 6 wishbone_out[24]
port 396 nsew signal output
rlabel metal2 s 71490 135200 71546 136000 6 wishbone_out[25]
port 397 nsew signal output
rlabel metal2 s 72226 135200 72282 136000 6 wishbone_out[26]
port 398 nsew signal output
rlabel metal2 s 73054 135200 73110 136000 6 wishbone_out[27]
port 399 nsew signal output
rlabel metal2 s 73882 135200 73938 136000 6 wishbone_out[28]
port 400 nsew signal output
rlabel metal2 s 74618 135200 74674 136000 6 wishbone_out[29]
port 401 nsew signal output
rlabel metal2 s 53366 135200 53422 136000 6 wishbone_out[2]
port 402 nsew signal output
rlabel metal2 s 75446 135200 75502 136000 6 wishbone_out[30]
port 403 nsew signal output
rlabel metal2 s 76182 135200 76238 136000 6 wishbone_out[31]
port 404 nsew signal output
rlabel metal2 s 77010 135200 77066 136000 6 wishbone_out[32]
port 405 nsew signal output
rlabel metal2 s 77746 135200 77802 136000 6 wishbone_out[33]
port 406 nsew signal output
rlabel metal2 s 78574 135200 78630 136000 6 wishbone_out[34]
port 407 nsew signal output
rlabel metal2 s 79310 135200 79366 136000 6 wishbone_out[35]
port 408 nsew signal output
rlabel metal2 s 80138 135200 80194 136000 6 wishbone_out[36]
port 409 nsew signal output
rlabel metal2 s 80874 135200 80930 136000 6 wishbone_out[37]
port 410 nsew signal output
rlabel metal2 s 81702 135200 81758 136000 6 wishbone_out[38]
port 411 nsew signal output
rlabel metal2 s 82530 135200 82586 136000 6 wishbone_out[39]
port 412 nsew signal output
rlabel metal2 s 54194 135200 54250 136000 6 wishbone_out[3]
port 413 nsew signal output
rlabel metal2 s 83266 135200 83322 136000 6 wishbone_out[40]
port 414 nsew signal output
rlabel metal2 s 84094 135200 84150 136000 6 wishbone_out[41]
port 415 nsew signal output
rlabel metal2 s 84830 135200 84886 136000 6 wishbone_out[42]
port 416 nsew signal output
rlabel metal2 s 85658 135200 85714 136000 6 wishbone_out[43]
port 417 nsew signal output
rlabel metal2 s 86394 135200 86450 136000 6 wishbone_out[44]
port 418 nsew signal output
rlabel metal2 s 87222 135200 87278 136000 6 wishbone_out[45]
port 419 nsew signal output
rlabel metal2 s 87958 135200 88014 136000 6 wishbone_out[46]
port 420 nsew signal output
rlabel metal2 s 88786 135200 88842 136000 6 wishbone_out[47]
port 421 nsew signal output
rlabel metal2 s 89522 135200 89578 136000 6 wishbone_out[48]
port 422 nsew signal output
rlabel metal2 s 90350 135200 90406 136000 6 wishbone_out[49]
port 423 nsew signal output
rlabel metal2 s 55022 135200 55078 136000 6 wishbone_out[4]
port 424 nsew signal output
rlabel metal2 s 91178 135200 91234 136000 6 wishbone_out[50]
port 425 nsew signal output
rlabel metal2 s 91914 135200 91970 136000 6 wishbone_out[51]
port 426 nsew signal output
rlabel metal2 s 92742 135200 92798 136000 6 wishbone_out[52]
port 427 nsew signal output
rlabel metal2 s 93478 135200 93534 136000 6 wishbone_out[53]
port 428 nsew signal output
rlabel metal2 s 94306 135200 94362 136000 6 wishbone_out[54]
port 429 nsew signal output
rlabel metal2 s 95042 135200 95098 136000 6 wishbone_out[55]
port 430 nsew signal output
rlabel metal2 s 95870 135200 95926 136000 6 wishbone_out[56]
port 431 nsew signal output
rlabel metal2 s 96606 135200 96662 136000 6 wishbone_out[57]
port 432 nsew signal output
rlabel metal2 s 97434 135200 97490 136000 6 wishbone_out[58]
port 433 nsew signal output
rlabel metal2 s 98170 135200 98226 136000 6 wishbone_out[59]
port 434 nsew signal output
rlabel metal2 s 55758 135200 55814 136000 6 wishbone_out[5]
port 435 nsew signal output
rlabel metal2 s 98998 135200 99054 136000 6 wishbone_out[60]
port 436 nsew signal output
rlabel metal2 s 99826 135200 99882 136000 6 wishbone_out[61]
port 437 nsew signal output
rlabel metal2 s 100562 135200 100618 136000 6 wishbone_out[62]
port 438 nsew signal output
rlabel metal2 s 101390 135200 101446 136000 6 wishbone_out[63]
port 439 nsew signal output
rlabel metal2 s 102126 135200 102182 136000 6 wishbone_out[64]
port 440 nsew signal output
rlabel metal2 s 102954 135200 103010 136000 6 wishbone_out[65]
port 441 nsew signal output
rlabel metal2 s 103690 135200 103746 136000 6 wishbone_out[66]
port 442 nsew signal output
rlabel metal2 s 104518 135200 104574 136000 6 wishbone_out[67]
port 443 nsew signal output
rlabel metal2 s 105254 135200 105310 136000 6 wishbone_out[68]
port 444 nsew signal output
rlabel metal2 s 106082 135200 106138 136000 6 wishbone_out[69]
port 445 nsew signal output
rlabel metal2 s 56586 135200 56642 136000 6 wishbone_out[6]
port 446 nsew signal output
rlabel metal2 s 106818 135200 106874 136000 6 wishbone_out[70]
port 447 nsew signal output
rlabel metal2 s 107646 135200 107702 136000 6 wishbone_out[71]
port 448 nsew signal output
rlabel metal2 s 108382 135200 108438 136000 6 wishbone_out[72]
port 449 nsew signal output
rlabel metal2 s 109210 135200 109266 136000 6 wishbone_out[73]
port 450 nsew signal output
rlabel metal2 s 110038 135200 110094 136000 6 wishbone_out[74]
port 451 nsew signal output
rlabel metal2 s 110774 135200 110830 136000 6 wishbone_out[75]
port 452 nsew signal output
rlabel metal2 s 111602 135200 111658 136000 6 wishbone_out[76]
port 453 nsew signal output
rlabel metal2 s 112338 135200 112394 136000 6 wishbone_out[77]
port 454 nsew signal output
rlabel metal2 s 113166 135200 113222 136000 6 wishbone_out[78]
port 455 nsew signal output
rlabel metal2 s 113902 135200 113958 136000 6 wishbone_out[79]
port 456 nsew signal output
rlabel metal2 s 57322 135200 57378 136000 6 wishbone_out[7]
port 457 nsew signal output
rlabel metal2 s 114730 135200 114786 136000 6 wishbone_out[80]
port 458 nsew signal output
rlabel metal2 s 115466 135200 115522 136000 6 wishbone_out[81]
port 459 nsew signal output
rlabel metal2 s 116294 135200 116350 136000 6 wishbone_out[82]
port 460 nsew signal output
rlabel metal2 s 117030 135200 117086 136000 6 wishbone_out[83]
port 461 nsew signal output
rlabel metal2 s 117858 135200 117914 136000 6 wishbone_out[84]
port 462 nsew signal output
rlabel metal2 s 118686 135200 118742 136000 6 wishbone_out[85]
port 463 nsew signal output
rlabel metal2 s 119422 135200 119478 136000 6 wishbone_out[86]
port 464 nsew signal output
rlabel metal2 s 120250 135200 120306 136000 6 wishbone_out[87]
port 465 nsew signal output
rlabel metal2 s 120986 135200 121042 136000 6 wishbone_out[88]
port 466 nsew signal output
rlabel metal2 s 121814 135200 121870 136000 6 wishbone_out[89]
port 467 nsew signal output
rlabel metal2 s 58150 135200 58206 136000 6 wishbone_out[8]
port 468 nsew signal output
rlabel metal2 s 122550 135200 122606 136000 6 wishbone_out[90]
port 469 nsew signal output
rlabel metal2 s 123378 135200 123434 136000 6 wishbone_out[91]
port 470 nsew signal output
rlabel metal2 s 124114 135200 124170 136000 6 wishbone_out[92]
port 471 nsew signal output
rlabel metal2 s 124942 135200 124998 136000 6 wishbone_out[93]
port 472 nsew signal output
rlabel metal2 s 125678 135200 125734 136000 6 wishbone_out[94]
port 473 nsew signal output
rlabel metal2 s 126506 135200 126562 136000 6 wishbone_out[95]
port 474 nsew signal output
rlabel metal2 s 127334 135200 127390 136000 6 wishbone_out[96]
port 475 nsew signal output
rlabel metal2 s 128070 135200 128126 136000 6 wishbone_out[97]
port 476 nsew signal output
rlabel metal2 s 128898 135200 128954 136000 6 wishbone_out[98]
port 477 nsew signal output
rlabel metal2 s 129634 135200 129690 136000 6 wishbone_out[99]
port 478 nsew signal output
rlabel metal2 s 58886 135200 58942 136000 6 wishbone_out[9]
port 479 nsew signal output
rlabel metal4 s 126708 2128 127028 133872 6 vccd1
port 480 nsew power bidirectional
rlabel metal4 s 95988 2128 96308 133872 6 vccd1
port 481 nsew power bidirectional
rlabel metal4 s 65268 2128 65588 133872 6 vccd1
port 482 nsew power bidirectional
rlabel metal4 s 34548 2128 34868 133872 6 vccd1
port 483 nsew power bidirectional
rlabel metal4 s 3828 2128 4148 133872 6 vccd1
port 484 nsew power bidirectional
rlabel metal4 s 111348 2128 111668 133872 6 vssd1
port 485 nsew ground bidirectional
rlabel metal4 s 80628 2128 80948 133872 6 vssd1
port 486 nsew ground bidirectional
rlabel metal4 s 49908 2128 50228 133872 6 vssd1
port 487 nsew ground bidirectional
rlabel metal4 s 19188 2128 19508 133872 6 vssd1
port 488 nsew ground bidirectional
rlabel metal4 s 127368 2176 127688 133824 6 vccd2
port 489 nsew power bidirectional
rlabel metal4 s 96648 2176 96968 133824 6 vccd2
port 490 nsew power bidirectional
rlabel metal4 s 65928 2176 66248 133824 6 vccd2
port 491 nsew power bidirectional
rlabel metal4 s 35208 2176 35528 133824 6 vccd2
port 492 nsew power bidirectional
rlabel metal4 s 4488 2176 4808 133824 6 vccd2
port 493 nsew power bidirectional
rlabel metal4 s 112008 2176 112328 133824 6 vssd2
port 494 nsew ground bidirectional
rlabel metal4 s 81288 2176 81608 133824 6 vssd2
port 495 nsew ground bidirectional
rlabel metal4 s 50568 2176 50888 133824 6 vssd2
port 496 nsew ground bidirectional
rlabel metal4 s 19848 2176 20168 133824 6 vssd2
port 497 nsew ground bidirectional
rlabel metal4 s 128028 2176 128348 133824 6 vdda1
port 498 nsew power bidirectional
rlabel metal4 s 97308 2176 97628 133824 6 vdda1
port 499 nsew power bidirectional
rlabel metal4 s 66588 2176 66908 133824 6 vdda1
port 500 nsew power bidirectional
rlabel metal4 s 35868 2176 36188 133824 6 vdda1
port 501 nsew power bidirectional
rlabel metal4 s 5148 2176 5468 133824 6 vdda1
port 502 nsew power bidirectional
rlabel metal4 s 112668 2176 112988 133824 6 vssa1
port 503 nsew ground bidirectional
rlabel metal4 s 81948 2176 82268 133824 6 vssa1
port 504 nsew ground bidirectional
rlabel metal4 s 51228 2176 51548 133824 6 vssa1
port 505 nsew ground bidirectional
rlabel metal4 s 20508 2176 20828 133824 6 vssa1
port 506 nsew ground bidirectional
rlabel metal4 s 128688 2176 129008 133824 6 vdda2
port 507 nsew power bidirectional
rlabel metal4 s 97968 2176 98288 133824 6 vdda2
port 508 nsew power bidirectional
rlabel metal4 s 67248 2176 67568 133824 6 vdda2
port 509 nsew power bidirectional
rlabel metal4 s 36528 2176 36848 133824 6 vdda2
port 510 nsew power bidirectional
rlabel metal4 s 5808 2176 6128 133824 6 vdda2
port 511 nsew power bidirectional
rlabel metal4 s 113328 2176 113648 133824 6 vssa2
port 512 nsew ground bidirectional
rlabel metal4 s 82608 2176 82928 133824 6 vssa2
port 513 nsew ground bidirectional
rlabel metal4 s 51888 2176 52208 133824 6 vssa2
port 514 nsew ground bidirectional
rlabel metal4 s 21168 2176 21488 133824 6 vssa2
port 515 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 1 0 135620 136000
string LEFview TRUE
string GDS_FILE /project/openlane/icache/runs/icache/results/magic/icache.gds
string GDS_END 50912432
string GDS_START 310896
<< end >>

