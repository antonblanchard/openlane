VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO multiply_4
  CLASS BLOCK ;
  FOREIGN multiply_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 798.550 BY 797.240 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.740 793.240 797.020 797.240 ;
    END
  END clk
  PIN m_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.020 793.240 0.300 797.240 ;
    END
  END m_in[0]
  PIN m_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.300 793.240 307.580 797.240 ;
    END
  END m_in[100]
  PIN m_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.520 793.240 310.800 797.240 ;
    END
  END m_in[101]
  PIN m_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.740 793.240 314.020 797.240 ;
    END
  END m_in[102]
  PIN m_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.500 793.240 316.780 797.240 ;
    END
  END m_in[103]
  PIN m_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.720 793.240 320.000 797.240 ;
    END
  END m_in[104]
  PIN m_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.940 793.240 323.220 797.240 ;
    END
  END m_in[105]
  PIN m_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.700 793.240 325.980 797.240 ;
    END
  END m_in[106]
  PIN m_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.920 793.240 329.200 797.240 ;
    END
  END m_in[107]
  PIN m_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.140 793.240 332.420 797.240 ;
    END
  END m_in[108]
  PIN m_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.360 793.240 335.640 797.240 ;
    END
  END m_in[109]
  PIN m_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.380 793.240 30.660 797.240 ;
    END
  END m_in[10]
  PIN m_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.120 793.240 338.400 797.240 ;
    END
  END m_in[110]
  PIN m_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.340 793.240 341.620 797.240 ;
    END
  END m_in[111]
  PIN m_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.560 793.240 344.840 797.240 ;
    END
  END m_in[112]
  PIN m_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.320 793.240 347.600 797.240 ;
    END
  END m_in[113]
  PIN m_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.540 793.240 350.820 797.240 ;
    END
  END m_in[114]
  PIN m_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.760 793.240 354.040 797.240 ;
    END
  END m_in[115]
  PIN m_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.520 793.240 356.800 797.240 ;
    END
  END m_in[116]
  PIN m_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.740 793.240 360.020 797.240 ;
    END
  END m_in[117]
  PIN m_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.960 793.240 363.240 797.240 ;
    END
  END m_in[118]
  PIN m_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.720 793.240 366.000 797.240 ;
    END
  END m_in[119]
  PIN m_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.600 793.240 33.880 797.240 ;
    END
  END m_in[11]
  PIN m_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.940 793.240 369.220 797.240 ;
    END
  END m_in[120]
  PIN m_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.160 793.240 372.440 797.240 ;
    END
  END m_in[121]
  PIN m_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.920 793.240 375.200 797.240 ;
    END
  END m_in[122]
  PIN m_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.140 793.240 378.420 797.240 ;
    END
  END m_in[123]
  PIN m_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.360 793.240 381.640 797.240 ;
    END
  END m_in[124]
  PIN m_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.580 793.240 384.860 797.240 ;
    END
  END m_in[125]
  PIN m_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.340 793.240 387.620 797.240 ;
    END
  END m_in[126]
  PIN m_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.560 793.240 390.840 797.240 ;
    END
  END m_in[127]
  PIN m_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.780 793.240 394.060 797.240 ;
    END
  END m_in[128]
  PIN m_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.540 793.240 396.820 797.240 ;
    END
  END m_in[129]
  PIN m_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.820 793.240 37.100 797.240 ;
    END
  END m_in[12]
  PIN m_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.760 793.240 400.040 797.240 ;
    END
  END m_in[130]
  PIN m_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.980 793.240 403.260 797.240 ;
    END
  END m_in[131]
  PIN m_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.740 793.240 406.020 797.240 ;
    END
  END m_in[132]
  PIN m_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.960 793.240 409.240 797.240 ;
    END
  END m_in[133]
  PIN m_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.180 793.240 412.460 797.240 ;
    END
  END m_in[134]
  PIN m_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.940 793.240 415.220 797.240 ;
    END
  END m_in[135]
  PIN m_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.160 793.240 418.440 797.240 ;
    END
  END m_in[136]
  PIN m_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.380 793.240 421.660 797.240 ;
    END
  END m_in[137]
  PIN m_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.600 793.240 424.880 797.240 ;
    END
  END m_in[138]
  PIN m_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.360 793.240 427.640 797.240 ;
    END
  END m_in[139]
  PIN m_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.580 793.240 39.860 797.240 ;
    END
  END m_in[13]
  PIN m_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.580 793.240 430.860 797.240 ;
    END
  END m_in[140]
  PIN m_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.800 793.240 434.080 797.240 ;
    END
  END m_in[141]
  PIN m_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.560 793.240 436.840 797.240 ;
    END
  END m_in[142]
  PIN m_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.780 793.240 440.060 797.240 ;
    END
  END m_in[143]
  PIN m_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.000 793.240 443.280 797.240 ;
    END
  END m_in[144]
  PIN m_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.760 793.240 446.040 797.240 ;
    END
  END m_in[145]
  PIN m_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.980 793.240 449.260 797.240 ;
    END
  END m_in[146]
  PIN m_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.200 793.240 452.480 797.240 ;
    END
  END m_in[147]
  PIN m_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.960 793.240 455.240 797.240 ;
    END
  END m_in[148]
  PIN m_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.180 793.240 458.460 797.240 ;
    END
  END m_in[149]
  PIN m_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.800 793.240 43.080 797.240 ;
    END
  END m_in[14]
  PIN m_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.400 793.240 461.680 797.240 ;
    END
  END m_in[150]
  PIN m_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.160 793.240 464.440 797.240 ;
    END
  END m_in[151]
  PIN m_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.380 793.240 467.660 797.240 ;
    END
  END m_in[152]
  PIN m_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.600 793.240 470.880 797.240 ;
    END
  END m_in[153]
  PIN m_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.820 793.240 474.100 797.240 ;
    END
  END m_in[154]
  PIN m_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.580 793.240 476.860 797.240 ;
    END
  END m_in[155]
  PIN m_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.800 793.240 480.080 797.240 ;
    END
  END m_in[156]
  PIN m_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.020 793.240 483.300 797.240 ;
    END
  END m_in[157]
  PIN m_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.780 793.240 486.060 797.240 ;
    END
  END m_in[158]
  PIN m_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.000 793.240 489.280 797.240 ;
    END
  END m_in[159]
  PIN m_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.020 793.240 46.300 797.240 ;
    END
  END m_in[15]
  PIN m_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.220 793.240 492.500 797.240 ;
    END
  END m_in[160]
  PIN m_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.980 793.240 495.260 797.240 ;
    END
  END m_in[161]
  PIN m_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.200 793.240 498.480 797.240 ;
    END
  END m_in[162]
  PIN m_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.420 793.240 501.700 797.240 ;
    END
  END m_in[163]
  PIN m_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.180 793.240 504.460 797.240 ;
    END
  END m_in[164]
  PIN m_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.400 793.240 507.680 797.240 ;
    END
  END m_in[165]
  PIN m_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.620 793.240 510.900 797.240 ;
    END
  END m_in[166]
  PIN m_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.380 793.240 513.660 797.240 ;
    END
  END m_in[167]
  PIN m_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.600 793.240 516.880 797.240 ;
    END
  END m_in[168]
  PIN m_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.820 793.240 520.100 797.240 ;
    END
  END m_in[169]
  PIN m_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.240 793.240 49.520 797.240 ;
    END
  END m_in[16]
  PIN m_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.040 793.240 523.320 797.240 ;
    END
  END m_in[170]
  PIN m_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.800 793.240 526.080 797.240 ;
    END
  END m_in[171]
  PIN m_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.020 793.240 529.300 797.240 ;
    END
  END m_in[172]
  PIN m_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.240 793.240 532.520 797.240 ;
    END
  END m_in[173]
  PIN m_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.000 793.240 535.280 797.240 ;
    END
  END m_in[174]
  PIN m_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.220 793.240 538.500 797.240 ;
    END
  END m_in[175]
  PIN m_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.440 793.240 541.720 797.240 ;
    END
  END m_in[176]
  PIN m_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.200 793.240 544.480 797.240 ;
    END
  END m_in[177]
  PIN m_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.420 793.240 547.700 797.240 ;
    END
  END m_in[178]
  PIN m_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.640 793.240 550.920 797.240 ;
    END
  END m_in[179]
  PIN m_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.000 793.240 52.280 797.240 ;
    END
  END m_in[17]
  PIN m_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.400 793.240 553.680 797.240 ;
    END
  END m_in[180]
  PIN m_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.620 793.240 556.900 797.240 ;
    END
  END m_in[181]
  PIN m_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.840 793.240 560.120 797.240 ;
    END
  END m_in[182]
  PIN m_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.600 793.240 562.880 797.240 ;
    END
  END m_in[183]
  PIN m_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.820 793.240 566.100 797.240 ;
    END
  END m_in[184]
  PIN m_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.040 793.240 569.320 797.240 ;
    END
  END m_in[185]
  PIN m_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.260 793.240 572.540 797.240 ;
    END
  END m_in[186]
  PIN m_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.020 793.240 575.300 797.240 ;
    END
  END m_in[187]
  PIN m_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.240 793.240 578.520 797.240 ;
    END
  END m_in[188]
  PIN m_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.460 793.240 581.740 797.240 ;
    END
  END m_in[189]
  PIN m_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.220 793.240 55.500 797.240 ;
    END
  END m_in[18]
  PIN m_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.220 793.240 584.500 797.240 ;
    END
  END m_in[190]
  PIN m_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.440 793.240 587.720 797.240 ;
    END
  END m_in[191]
  PIN m_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.660 793.240 590.940 797.240 ;
    END
  END m_in[192]
  PIN m_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.420 793.240 593.700 797.240 ;
    END
  END m_in[193]
  PIN m_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.640 793.240 596.920 797.240 ;
    END
  END m_in[194]
  PIN m_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.860 793.240 600.140 797.240 ;
    END
  END m_in[195]
  PIN m_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.620 793.240 602.900 797.240 ;
    END
  END m_in[196]
  PIN m_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.840 793.240 606.120 797.240 ;
    END
  END m_in[197]
  PIN m_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.060 793.240 609.340 797.240 ;
    END
  END m_in[198]
  PIN m_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.280 793.240 612.560 797.240 ;
    END
  END m_in[199]
  PIN m_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.440 793.240 58.720 797.240 ;
    END
  END m_in[19]
  PIN m_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.780 793.240 3.060 797.240 ;
    END
  END m_in[1]
  PIN m_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.040 793.240 615.320 797.240 ;
    END
  END m_in[200]
  PIN m_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.260 793.240 618.540 797.240 ;
    END
  END m_in[201]
  PIN m_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.480 793.240 621.760 797.240 ;
    END
  END m_in[202]
  PIN m_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.240 793.240 624.520 797.240 ;
    END
  END m_in[203]
  PIN m_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.460 793.240 627.740 797.240 ;
    END
  END m_in[204]
  PIN m_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.680 793.240 630.960 797.240 ;
    END
  END m_in[205]
  PIN m_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.440 793.240 633.720 797.240 ;
    END
  END m_in[206]
  PIN m_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.660 793.240 636.940 797.240 ;
    END
  END m_in[207]
  PIN m_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.880 793.240 640.160 797.240 ;
    END
  END m_in[208]
  PIN m_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.640 793.240 642.920 797.240 ;
    END
  END m_in[209]
  PIN m_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.200 793.240 61.480 797.240 ;
    END
  END m_in[20]
  PIN m_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.860 793.240 646.140 797.240 ;
    END
  END m_in[210]
  PIN m_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.080 793.240 649.360 797.240 ;
    END
  END m_in[211]
  PIN m_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.840 793.240 652.120 797.240 ;
    END
  END m_in[212]
  PIN m_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.060 793.240 655.340 797.240 ;
    END
  END m_in[213]
  PIN m_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.280 793.240 658.560 797.240 ;
    END
  END m_in[214]
  PIN m_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.500 793.240 661.780 797.240 ;
    END
  END m_in[215]
  PIN m_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.260 793.240 664.540 797.240 ;
    END
  END m_in[216]
  PIN m_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.480 793.240 667.760 797.240 ;
    END
  END m_in[217]
  PIN m_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.700 793.240 670.980 797.240 ;
    END
  END m_in[218]
  PIN m_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.460 793.240 673.740 797.240 ;
    END
  END m_in[219]
  PIN m_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.420 793.240 64.700 797.240 ;
    END
  END m_in[21]
  PIN m_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.680 793.240 676.960 797.240 ;
    END
  END m_in[220]
  PIN m_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.900 793.240 680.180 797.240 ;
    END
  END m_in[221]
  PIN m_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.660 793.240 682.940 797.240 ;
    END
  END m_in[222]
  PIN m_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.880 793.240 686.160 797.240 ;
    END
  END m_in[223]
  PIN m_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.100 793.240 689.380 797.240 ;
    END
  END m_in[224]
  PIN m_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.860 793.240 692.140 797.240 ;
    END
  END m_in[225]
  PIN m_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.080 793.240 695.360 797.240 ;
    END
  END m_in[226]
  PIN m_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.300 793.240 698.580 797.240 ;
    END
  END m_in[227]
  PIN m_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.060 793.240 701.340 797.240 ;
    END
  END m_in[228]
  PIN m_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.280 793.240 704.560 797.240 ;
    END
  END m_in[229]
  PIN m_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.640 793.240 67.920 797.240 ;
    END
  END m_in[22]
  PIN m_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.500 793.240 707.780 797.240 ;
    END
  END m_in[230]
  PIN m_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.720 793.240 711.000 797.240 ;
    END
  END m_in[231]
  PIN m_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.480 793.240 713.760 797.240 ;
    END
  END m_in[232]
  PIN m_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.700 793.240 716.980 797.240 ;
    END
  END m_in[233]
  PIN m_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.920 793.240 720.200 797.240 ;
    END
  END m_in[234]
  PIN m_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.680 793.240 722.960 797.240 ;
    END
  END m_in[235]
  PIN m_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.900 793.240 726.180 797.240 ;
    END
  END m_in[236]
  PIN m_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.120 793.240 729.400 797.240 ;
    END
  END m_in[237]
  PIN m_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.880 793.240 732.160 797.240 ;
    END
  END m_in[238]
  PIN m_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.100 793.240 735.380 797.240 ;
    END
  END m_in[239]
  PIN m_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.400 793.240 70.680 797.240 ;
    END
  END m_in[23]
  PIN m_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.320 793.240 738.600 797.240 ;
    END
  END m_in[240]
  PIN m_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.080 793.240 741.360 797.240 ;
    END
  END m_in[241]
  PIN m_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.300 793.240 744.580 797.240 ;
    END
  END m_in[242]
  PIN m_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.520 793.240 747.800 797.240 ;
    END
  END m_in[243]
  PIN m_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.280 793.240 750.560 797.240 ;
    END
  END m_in[244]
  PIN m_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.500 793.240 753.780 797.240 ;
    END
  END m_in[245]
  PIN m_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.720 793.240 757.000 797.240 ;
    END
  END m_in[246]
  PIN m_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.940 793.240 760.220 797.240 ;
    END
  END m_in[247]
  PIN m_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.700 793.240 762.980 797.240 ;
    END
  END m_in[248]
  PIN m_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.920 793.240 766.200 797.240 ;
    END
  END m_in[249]
  PIN m_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.620 793.240 73.900 797.240 ;
    END
  END m_in[24]
  PIN m_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.140 793.240 769.420 797.240 ;
    END
  END m_in[250]
  PIN m_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.900 793.240 772.180 797.240 ;
    END
  END m_in[251]
  PIN m_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.120 793.240 775.400 797.240 ;
    END
  END m_in[252]
  PIN m_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.340 793.240 778.620 797.240 ;
    END
  END m_in[253]
  PIN m_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.100 793.240 781.380 797.240 ;
    END
  END m_in[254]
  PIN m_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.320 793.240 784.600 797.240 ;
    END
  END m_in[255]
  PIN m_in[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.540 793.240 787.820 797.240 ;
    END
  END m_in[256]
  PIN m_in[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.300 793.240 790.580 797.240 ;
    END
  END m_in[257]
  PIN m_in[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.520 793.240 793.800 797.240 ;
    END
  END m_in[258]
  PIN m_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.840 793.240 77.120 797.240 ;
    END
  END m_in[25]
  PIN m_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.600 793.240 79.880 797.240 ;
    END
  END m_in[26]
  PIN m_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.820 793.240 83.100 797.240 ;
    END
  END m_in[27]
  PIN m_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.040 793.240 86.320 797.240 ;
    END
  END m_in[28]
  PIN m_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.800 793.240 89.080 797.240 ;
    END
  END m_in[29]
  PIN m_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.000 793.240 6.280 797.240 ;
    END
  END m_in[2]
  PIN m_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.020 793.240 92.300 797.240 ;
    END
  END m_in[30]
  PIN m_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.240 793.240 95.520 797.240 ;
    END
  END m_in[31]
  PIN m_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.460 793.240 98.740 797.240 ;
    END
  END m_in[32]
  PIN m_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.220 793.240 101.500 797.240 ;
    END
  END m_in[33]
  PIN m_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.440 793.240 104.720 797.240 ;
    END
  END m_in[34]
  PIN m_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.660 793.240 107.940 797.240 ;
    END
  END m_in[35]
  PIN m_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.420 793.240 110.700 797.240 ;
    END
  END m_in[36]
  PIN m_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.640 793.240 113.920 797.240 ;
    END
  END m_in[37]
  PIN m_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.860 793.240 117.140 797.240 ;
    END
  END m_in[38]
  PIN m_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.620 793.240 119.900 797.240 ;
    END
  END m_in[39]
  PIN m_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.220 793.240 9.500 797.240 ;
    END
  END m_in[3]
  PIN m_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.840 793.240 123.120 797.240 ;
    END
  END m_in[40]
  PIN m_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.060 793.240 126.340 797.240 ;
    END
  END m_in[41]
  PIN m_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.820 793.240 129.100 797.240 ;
    END
  END m_in[42]
  PIN m_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.040 793.240 132.320 797.240 ;
    END
  END m_in[43]
  PIN m_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.260 793.240 135.540 797.240 ;
    END
  END m_in[44]
  PIN m_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.020 793.240 138.300 797.240 ;
    END
  END m_in[45]
  PIN m_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.240 793.240 141.520 797.240 ;
    END
  END m_in[46]
  PIN m_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.460 793.240 144.740 797.240 ;
    END
  END m_in[47]
  PIN m_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.680 793.240 147.960 797.240 ;
    END
  END m_in[48]
  PIN m_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.440 793.240 150.720 797.240 ;
    END
  END m_in[49]
  PIN m_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.980 793.240 12.260 797.240 ;
    END
  END m_in[4]
  PIN m_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.660 793.240 153.940 797.240 ;
    END
  END m_in[50]
  PIN m_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.880 793.240 157.160 797.240 ;
    END
  END m_in[51]
  PIN m_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.640 793.240 159.920 797.240 ;
    END
  END m_in[52]
  PIN m_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.860 793.240 163.140 797.240 ;
    END
  END m_in[53]
  PIN m_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.080 793.240 166.360 797.240 ;
    END
  END m_in[54]
  PIN m_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.840 793.240 169.120 797.240 ;
    END
  END m_in[55]
  PIN m_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.060 793.240 172.340 797.240 ;
    END
  END m_in[56]
  PIN m_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.280 793.240 175.560 797.240 ;
    END
  END m_in[57]
  PIN m_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.040 793.240 178.320 797.240 ;
    END
  END m_in[58]
  PIN m_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.260 793.240 181.540 797.240 ;
    END
  END m_in[59]
  PIN m_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.200 793.240 15.480 797.240 ;
    END
  END m_in[5]
  PIN m_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.480 793.240 184.760 797.240 ;
    END
  END m_in[60]
  PIN m_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.240 793.240 187.520 797.240 ;
    END
  END m_in[61]
  PIN m_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.460 793.240 190.740 797.240 ;
    END
  END m_in[62]
  PIN m_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.680 793.240 193.960 797.240 ;
    END
  END m_in[63]
  PIN m_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.900 793.240 197.180 797.240 ;
    END
  END m_in[64]
  PIN m_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.660 793.240 199.940 797.240 ;
    END
  END m_in[65]
  PIN m_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.880 793.240 203.160 797.240 ;
    END
  END m_in[66]
  PIN m_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.100 793.240 206.380 797.240 ;
    END
  END m_in[67]
  PIN m_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.860 793.240 209.140 797.240 ;
    END
  END m_in[68]
  PIN m_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.080 793.240 212.360 797.240 ;
    END
  END m_in[69]
  PIN m_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.420 793.240 18.700 797.240 ;
    END
  END m_in[6]
  PIN m_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.300 793.240 215.580 797.240 ;
    END
  END m_in[70]
  PIN m_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.060 793.240 218.340 797.240 ;
    END
  END m_in[71]
  PIN m_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.280 793.240 221.560 797.240 ;
    END
  END m_in[72]
  PIN m_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.500 793.240 224.780 797.240 ;
    END
  END m_in[73]
  PIN m_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.260 793.240 227.540 797.240 ;
    END
  END m_in[74]
  PIN m_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.480 793.240 230.760 797.240 ;
    END
  END m_in[75]
  PIN m_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.700 793.240 233.980 797.240 ;
    END
  END m_in[76]
  PIN m_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.920 793.240 237.200 797.240 ;
    END
  END m_in[77]
  PIN m_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.680 793.240 239.960 797.240 ;
    END
  END m_in[78]
  PIN m_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.900 793.240 243.180 797.240 ;
    END
  END m_in[79]
  PIN m_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.180 793.240 21.460 797.240 ;
    END
  END m_in[7]
  PIN m_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.120 793.240 246.400 797.240 ;
    END
  END m_in[80]
  PIN m_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.880 793.240 249.160 797.240 ;
    END
  END m_in[81]
  PIN m_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.100 793.240 252.380 797.240 ;
    END
  END m_in[82]
  PIN m_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.320 793.240 255.600 797.240 ;
    END
  END m_in[83]
  PIN m_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.080 793.240 258.360 797.240 ;
    END
  END m_in[84]
  PIN m_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.300 793.240 261.580 797.240 ;
    END
  END m_in[85]
  PIN m_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.520 793.240 264.800 797.240 ;
    END
  END m_in[86]
  PIN m_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.280 793.240 267.560 797.240 ;
    END
  END m_in[87]
  PIN m_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.500 793.240 270.780 797.240 ;
    END
  END m_in[88]
  PIN m_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.720 793.240 274.000 797.240 ;
    END
  END m_in[89]
  PIN m_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.400 793.240 24.680 797.240 ;
    END
  END m_in[8]
  PIN m_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.480 793.240 276.760 797.240 ;
    END
  END m_in[90]
  PIN m_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.700 793.240 279.980 797.240 ;
    END
  END m_in[91]
  PIN m_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.920 793.240 283.200 797.240 ;
    END
  END m_in[92]
  PIN m_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.140 793.240 286.420 797.240 ;
    END
  END m_in[93]
  PIN m_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.900 793.240 289.180 797.240 ;
    END
  END m_in[94]
  PIN m_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.120 793.240 292.400 797.240 ;
    END
  END m_in[95]
  PIN m_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.340 793.240 295.620 797.240 ;
    END
  END m_in[96]
  PIN m_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.100 793.240 298.380 797.240 ;
    END
  END m_in[97]
  PIN m_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.320 793.240 301.600 797.240 ;
    END
  END m_in[98]
  PIN m_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.540 793.240 304.820 797.240 ;
    END
  END m_in[99]
  PIN m_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.620 793.240 27.900 797.240 ;
    END
  END m_in[9]
  PIN m_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 0.000 798.550 0.600 ;
    END
  END m_out[0]
  PIN m_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 614.720 798.550 615.320 ;
    END
  END m_out[100]
  PIN m_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 620.840 798.550 621.440 ;
    END
  END m_out[101]
  PIN m_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 626.960 798.550 627.560 ;
    END
  END m_out[102]
  PIN m_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 633.080 798.550 633.680 ;
    END
  END m_out[103]
  PIN m_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 639.200 798.550 639.800 ;
    END
  END m_out[104]
  PIN m_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 645.320 798.550 645.920 ;
    END
  END m_out[105]
  PIN m_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 651.440 798.550 652.040 ;
    END
  END m_out[106]
  PIN m_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 657.560 798.550 658.160 ;
    END
  END m_out[107]
  PIN m_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 663.680 798.550 664.280 ;
    END
  END m_out[108]
  PIN m_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 670.480 798.550 671.080 ;
    END
  END m_out[109]
  PIN m_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 61.200 798.550 61.800 ;
    END
  END m_out[10]
  PIN m_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 676.600 798.550 677.200 ;
    END
  END m_out[110]
  PIN m_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 682.720 798.550 683.320 ;
    END
  END m_out[111]
  PIN m_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 688.840 798.550 689.440 ;
    END
  END m_out[112]
  PIN m_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 694.960 798.550 695.560 ;
    END
  END m_out[113]
  PIN m_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 701.080 798.550 701.680 ;
    END
  END m_out[114]
  PIN m_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 707.200 798.550 707.800 ;
    END
  END m_out[115]
  PIN m_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 713.320 798.550 713.920 ;
    END
  END m_out[116]
  PIN m_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 719.440 798.550 720.040 ;
    END
  END m_out[117]
  PIN m_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 725.560 798.550 726.160 ;
    END
  END m_out[118]
  PIN m_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 731.680 798.550 732.280 ;
    END
  END m_out[119]
  PIN m_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 67.320 798.550 67.920 ;
    END
  END m_out[11]
  PIN m_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 737.800 798.550 738.400 ;
    END
  END m_out[120]
  PIN m_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 743.920 798.550 744.520 ;
    END
  END m_out[121]
  PIN m_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 750.040 798.550 750.640 ;
    END
  END m_out[122]
  PIN m_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 756.160 798.550 756.760 ;
    END
  END m_out[123]
  PIN m_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 762.280 798.550 762.880 ;
    END
  END m_out[124]
  PIN m_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 768.400 798.550 769.000 ;
    END
  END m_out[125]
  PIN m_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 774.520 798.550 775.120 ;
    END
  END m_out[126]
  PIN m_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 780.640 798.550 781.240 ;
    END
  END m_out[127]
  PIN m_out[128]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 786.760 798.550 787.360 ;
    END
  END m_out[128]
  PIN m_out[129]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 792.880 798.550 793.480 ;
    END
  END m_out[129]
  PIN m_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 73.440 798.550 74.040 ;
    END
  END m_out[12]
  PIN m_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 79.560 798.550 80.160 ;
    END
  END m_out[13]
  PIN m_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 85.680 798.550 86.280 ;
    END
  END m_out[14]
  PIN m_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 91.800 798.550 92.400 ;
    END
  END m_out[15]
  PIN m_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 97.920 798.550 98.520 ;
    END
  END m_out[16]
  PIN m_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 104.040 798.550 104.640 ;
    END
  END m_out[17]
  PIN m_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 110.160 798.550 110.760 ;
    END
  END m_out[18]
  PIN m_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 116.280 798.550 116.880 ;
    END
  END m_out[19]
  PIN m_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 6.120 798.550 6.720 ;
    END
  END m_out[1]
  PIN m_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 122.400 798.550 123.000 ;
    END
  END m_out[20]
  PIN m_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 128.520 798.550 129.120 ;
    END
  END m_out[21]
  PIN m_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 135.320 798.550 135.920 ;
    END
  END m_out[22]
  PIN m_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 141.440 798.550 142.040 ;
    END
  END m_out[23]
  PIN m_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 147.560 798.550 148.160 ;
    END
  END m_out[24]
  PIN m_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 153.680 798.550 154.280 ;
    END
  END m_out[25]
  PIN m_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 159.800 798.550 160.400 ;
    END
  END m_out[26]
  PIN m_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 165.920 798.550 166.520 ;
    END
  END m_out[27]
  PIN m_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 172.040 798.550 172.640 ;
    END
  END m_out[28]
  PIN m_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 178.160 798.550 178.760 ;
    END
  END m_out[29]
  PIN m_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 12.240 798.550 12.840 ;
    END
  END m_out[2]
  PIN m_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 184.280 798.550 184.880 ;
    END
  END m_out[30]
  PIN m_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 190.400 798.550 191.000 ;
    END
  END m_out[31]
  PIN m_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 196.520 798.550 197.120 ;
    END
  END m_out[32]
  PIN m_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 202.640 798.550 203.240 ;
    END
  END m_out[33]
  PIN m_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 208.760 798.550 209.360 ;
    END
  END m_out[34]
  PIN m_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 214.880 798.550 215.480 ;
    END
  END m_out[35]
  PIN m_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 221.000 798.550 221.600 ;
    END
  END m_out[36]
  PIN m_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 227.120 798.550 227.720 ;
    END
  END m_out[37]
  PIN m_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 233.240 798.550 233.840 ;
    END
  END m_out[38]
  PIN m_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 239.360 798.550 239.960 ;
    END
  END m_out[39]
  PIN m_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 18.360 798.550 18.960 ;
    END
  END m_out[3]
  PIN m_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 245.480 798.550 246.080 ;
    END
  END m_out[40]
  PIN m_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 251.600 798.550 252.200 ;
    END
  END m_out[41]
  PIN m_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 257.720 798.550 258.320 ;
    END
  END m_out[42]
  PIN m_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 263.840 798.550 264.440 ;
    END
  END m_out[43]
  PIN m_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 270.640 798.550 271.240 ;
    END
  END m_out[44]
  PIN m_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 276.760 798.550 277.360 ;
    END
  END m_out[45]
  PIN m_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 282.880 798.550 283.480 ;
    END
  END m_out[46]
  PIN m_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 289.000 798.550 289.600 ;
    END
  END m_out[47]
  PIN m_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 295.120 798.550 295.720 ;
    END
  END m_out[48]
  PIN m_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 301.240 798.550 301.840 ;
    END
  END m_out[49]
  PIN m_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 24.480 798.550 25.080 ;
    END
  END m_out[4]
  PIN m_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 307.360 798.550 307.960 ;
    END
  END m_out[50]
  PIN m_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 313.480 798.550 314.080 ;
    END
  END m_out[51]
  PIN m_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 319.600 798.550 320.200 ;
    END
  END m_out[52]
  PIN m_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 325.720 798.550 326.320 ;
    END
  END m_out[53]
  PIN m_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 331.840 798.550 332.440 ;
    END
  END m_out[54]
  PIN m_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 337.960 798.550 338.560 ;
    END
  END m_out[55]
  PIN m_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 344.080 798.550 344.680 ;
    END
  END m_out[56]
  PIN m_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 350.200 798.550 350.800 ;
    END
  END m_out[57]
  PIN m_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 356.320 798.550 356.920 ;
    END
  END m_out[58]
  PIN m_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 362.440 798.550 363.040 ;
    END
  END m_out[59]
  PIN m_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 30.600 798.550 31.200 ;
    END
  END m_out[5]
  PIN m_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 368.560 798.550 369.160 ;
    END
  END m_out[60]
  PIN m_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 374.680 798.550 375.280 ;
    END
  END m_out[61]
  PIN m_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 380.800 798.550 381.400 ;
    END
  END m_out[62]
  PIN m_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 386.920 798.550 387.520 ;
    END
  END m_out[63]
  PIN m_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 393.040 798.550 393.640 ;
    END
  END m_out[64]
  PIN m_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 399.840 798.550 400.440 ;
    END
  END m_out[65]
  PIN m_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 405.960 798.550 406.560 ;
    END
  END m_out[66]
  PIN m_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 412.080 798.550 412.680 ;
    END
  END m_out[67]
  PIN m_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 418.200 798.550 418.800 ;
    END
  END m_out[68]
  PIN m_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 424.320 798.550 424.920 ;
    END
  END m_out[69]
  PIN m_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 36.720 798.550 37.320 ;
    END
  END m_out[6]
  PIN m_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 430.440 798.550 431.040 ;
    END
  END m_out[70]
  PIN m_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 436.560 798.550 437.160 ;
    END
  END m_out[71]
  PIN m_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 442.680 798.550 443.280 ;
    END
  END m_out[72]
  PIN m_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 448.800 798.550 449.400 ;
    END
  END m_out[73]
  PIN m_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 454.920 798.550 455.520 ;
    END
  END m_out[74]
  PIN m_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 461.040 798.550 461.640 ;
    END
  END m_out[75]
  PIN m_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 467.160 798.550 467.760 ;
    END
  END m_out[76]
  PIN m_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 473.280 798.550 473.880 ;
    END
  END m_out[77]
  PIN m_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 479.400 798.550 480.000 ;
    END
  END m_out[78]
  PIN m_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 485.520 798.550 486.120 ;
    END
  END m_out[79]
  PIN m_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 42.840 798.550 43.440 ;
    END
  END m_out[7]
  PIN m_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 491.640 798.550 492.240 ;
    END
  END m_out[80]
  PIN m_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 497.760 798.550 498.360 ;
    END
  END m_out[81]
  PIN m_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 503.880 798.550 504.480 ;
    END
  END m_out[82]
  PIN m_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 510.000 798.550 510.600 ;
    END
  END m_out[83]
  PIN m_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 516.120 798.550 516.720 ;
    END
  END m_out[84]
  PIN m_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 522.240 798.550 522.840 ;
    END
  END m_out[85]
  PIN m_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 528.360 798.550 528.960 ;
    END
  END m_out[86]
  PIN m_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 535.160 798.550 535.760 ;
    END
  END m_out[87]
  PIN m_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 541.280 798.550 541.880 ;
    END
  END m_out[88]
  PIN m_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 547.400 798.550 548.000 ;
    END
  END m_out[89]
  PIN m_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 48.960 798.550 49.560 ;
    END
  END m_out[8]
  PIN m_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 553.520 798.550 554.120 ;
    END
  END m_out[90]
  PIN m_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 559.640 798.550 560.240 ;
    END
  END m_out[91]
  PIN m_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 565.760 798.550 566.360 ;
    END
  END m_out[92]
  PIN m_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 571.880 798.550 572.480 ;
    END
  END m_out[93]
  PIN m_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 578.000 798.550 578.600 ;
    END
  END m_out[94]
  PIN m_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 584.120 798.550 584.720 ;
    END
  END m_out[95]
  PIN m_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 590.240 798.550 590.840 ;
    END
  END m_out[96]
  PIN m_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 596.360 798.550 596.960 ;
    END
  END m_out[97]
  PIN m_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 602.480 798.550 603.080 ;
    END
  END m_out[98]
  PIN m_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 608.600 798.550 609.200 ;
    END
  END m_out[99]
  PIN m_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.550 55.080 798.550 55.680 ;
    END
  END m_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 787.590 7.880 789.190 786.280 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 633.990 7.880 635.590 786.280 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 480.390 7.880 481.990 786.280 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 326.790 7.880 328.390 786.280 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 173.190 7.880 174.790 786.280 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.590 7.880 21.190 786.280 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 710.790 7.880 712.390 786.280 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 557.190 7.880 558.790 786.280 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 403.590 7.880 405.190 786.280 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 249.990 7.880 251.590 786.280 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.390 7.880 97.990 786.280 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 637.290 8.120 638.890 786.040 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 483.690 8.120 485.290 786.040 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 330.090 8.120 331.690 786.040 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 176.490 8.120 178.090 786.040 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.890 8.120 24.490 786.040 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 714.090 8.120 715.690 786.040 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 560.490 8.120 562.090 786.040 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 406.890 8.120 408.490 786.040 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 253.290 8.120 254.890 786.040 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 99.690 8.120 101.290 786.040 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 640.590 8.120 642.190 786.040 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 486.990 8.120 488.590 786.040 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 333.390 8.120 334.990 786.040 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 179.790 8.120 181.390 786.040 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 26.190 8.120 27.790 786.040 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 717.390 8.120 718.990 786.040 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 563.790 8.120 565.390 786.040 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 410.190 8.120 411.790 786.040 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 256.590 8.120 258.190 786.040 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 102.990 8.120 104.590 786.040 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 643.890 8.120 645.490 786.040 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 490.290 8.120 491.890 786.040 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 336.690 8.120 338.290 786.040 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 183.090 8.120 184.690 786.040 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 29.490 8.120 31.090 786.040 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 720.690 8.120 722.290 786.040 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 567.090 8.120 568.690 786.040 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 413.490 8.120 415.090 786.040 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 259.890 8.120 261.490 786.040 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 106.290 8.120 107.890 786.040 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 4.070 8.035 793.745 791.395 ;
      LAYER met1 ;
        RECT 0.000 5.440 797.040 791.440 ;
      LAYER met2 ;
        RECT 0.580 792.960 2.500 793.365 ;
        RECT 3.340 792.960 5.720 793.365 ;
        RECT 6.560 792.960 8.940 793.365 ;
        RECT 9.780 792.960 11.700 793.365 ;
        RECT 12.540 792.960 14.920 793.365 ;
        RECT 15.760 792.960 18.140 793.365 ;
        RECT 18.980 792.960 20.900 793.365 ;
        RECT 21.740 792.960 24.120 793.365 ;
        RECT 24.960 792.960 27.340 793.365 ;
        RECT 28.180 792.960 30.100 793.365 ;
        RECT 30.940 792.960 33.320 793.365 ;
        RECT 34.160 792.960 36.540 793.365 ;
        RECT 37.380 792.960 39.300 793.365 ;
        RECT 40.140 792.960 42.520 793.365 ;
        RECT 43.360 792.960 45.740 793.365 ;
        RECT 46.580 792.960 48.960 793.365 ;
        RECT 49.800 792.960 51.720 793.365 ;
        RECT 52.560 792.960 54.940 793.365 ;
        RECT 55.780 792.960 58.160 793.365 ;
        RECT 59.000 792.960 60.920 793.365 ;
        RECT 61.760 792.960 64.140 793.365 ;
        RECT 64.980 792.960 67.360 793.365 ;
        RECT 68.200 792.960 70.120 793.365 ;
        RECT 70.960 792.960 73.340 793.365 ;
        RECT 74.180 792.960 76.560 793.365 ;
        RECT 77.400 792.960 79.320 793.365 ;
        RECT 80.160 792.960 82.540 793.365 ;
        RECT 83.380 792.960 85.760 793.365 ;
        RECT 86.600 792.960 88.520 793.365 ;
        RECT 89.360 792.960 91.740 793.365 ;
        RECT 92.580 792.960 94.960 793.365 ;
        RECT 95.800 792.960 98.180 793.365 ;
        RECT 99.020 792.960 100.940 793.365 ;
        RECT 101.780 792.960 104.160 793.365 ;
        RECT 105.000 792.960 107.380 793.365 ;
        RECT 108.220 792.960 110.140 793.365 ;
        RECT 110.980 792.960 113.360 793.365 ;
        RECT 114.200 792.960 116.580 793.365 ;
        RECT 117.420 792.960 119.340 793.365 ;
        RECT 120.180 792.960 122.560 793.365 ;
        RECT 123.400 792.960 125.780 793.365 ;
        RECT 126.620 792.960 128.540 793.365 ;
        RECT 129.380 792.960 131.760 793.365 ;
        RECT 132.600 792.960 134.980 793.365 ;
        RECT 135.820 792.960 137.740 793.365 ;
        RECT 138.580 792.960 140.960 793.365 ;
        RECT 141.800 792.960 144.180 793.365 ;
        RECT 145.020 792.960 147.400 793.365 ;
        RECT 148.240 792.960 150.160 793.365 ;
        RECT 151.000 792.960 153.380 793.365 ;
        RECT 154.220 792.960 156.600 793.365 ;
        RECT 157.440 792.960 159.360 793.365 ;
        RECT 160.200 792.960 162.580 793.365 ;
        RECT 163.420 792.960 165.800 793.365 ;
        RECT 166.640 792.960 168.560 793.365 ;
        RECT 169.400 792.960 171.780 793.365 ;
        RECT 172.620 792.960 175.000 793.365 ;
        RECT 175.840 792.960 177.760 793.365 ;
        RECT 178.600 792.960 180.980 793.365 ;
        RECT 181.820 792.960 184.200 793.365 ;
        RECT 185.040 792.960 186.960 793.365 ;
        RECT 187.800 792.960 190.180 793.365 ;
        RECT 191.020 792.960 193.400 793.365 ;
        RECT 194.240 792.960 196.620 793.365 ;
        RECT 197.460 792.960 199.380 793.365 ;
        RECT 200.220 792.960 202.600 793.365 ;
        RECT 203.440 792.960 205.820 793.365 ;
        RECT 206.660 792.960 208.580 793.365 ;
        RECT 209.420 792.960 211.800 793.365 ;
        RECT 212.640 792.960 215.020 793.365 ;
        RECT 215.860 792.960 217.780 793.365 ;
        RECT 218.620 792.960 221.000 793.365 ;
        RECT 221.840 792.960 224.220 793.365 ;
        RECT 225.060 792.960 226.980 793.365 ;
        RECT 227.820 792.960 230.200 793.365 ;
        RECT 231.040 792.960 233.420 793.365 ;
        RECT 234.260 792.960 236.640 793.365 ;
        RECT 237.480 792.960 239.400 793.365 ;
        RECT 240.240 792.960 242.620 793.365 ;
        RECT 243.460 792.960 245.840 793.365 ;
        RECT 246.680 792.960 248.600 793.365 ;
        RECT 249.440 792.960 251.820 793.365 ;
        RECT 252.660 792.960 255.040 793.365 ;
        RECT 255.880 792.960 257.800 793.365 ;
        RECT 258.640 792.960 261.020 793.365 ;
        RECT 261.860 792.960 264.240 793.365 ;
        RECT 265.080 792.960 267.000 793.365 ;
        RECT 267.840 792.960 270.220 793.365 ;
        RECT 271.060 792.960 273.440 793.365 ;
        RECT 274.280 792.960 276.200 793.365 ;
        RECT 277.040 792.960 279.420 793.365 ;
        RECT 280.260 792.960 282.640 793.365 ;
        RECT 283.480 792.960 285.860 793.365 ;
        RECT 286.700 792.960 288.620 793.365 ;
        RECT 289.460 792.960 291.840 793.365 ;
        RECT 292.680 792.960 295.060 793.365 ;
        RECT 295.900 792.960 297.820 793.365 ;
        RECT 298.660 792.960 301.040 793.365 ;
        RECT 301.880 792.960 304.260 793.365 ;
        RECT 305.100 792.960 307.020 793.365 ;
        RECT 307.860 792.960 310.240 793.365 ;
        RECT 311.080 792.960 313.460 793.365 ;
        RECT 314.300 792.960 316.220 793.365 ;
        RECT 317.060 792.960 319.440 793.365 ;
        RECT 320.280 792.960 322.660 793.365 ;
        RECT 323.500 792.960 325.420 793.365 ;
        RECT 326.260 792.960 328.640 793.365 ;
        RECT 329.480 792.960 331.860 793.365 ;
        RECT 332.700 792.960 335.080 793.365 ;
        RECT 335.920 792.960 337.840 793.365 ;
        RECT 338.680 792.960 341.060 793.365 ;
        RECT 341.900 792.960 344.280 793.365 ;
        RECT 345.120 792.960 347.040 793.365 ;
        RECT 347.880 792.960 350.260 793.365 ;
        RECT 351.100 792.960 353.480 793.365 ;
        RECT 354.320 792.960 356.240 793.365 ;
        RECT 357.080 792.960 359.460 793.365 ;
        RECT 360.300 792.960 362.680 793.365 ;
        RECT 363.520 792.960 365.440 793.365 ;
        RECT 366.280 792.960 368.660 793.365 ;
        RECT 369.500 792.960 371.880 793.365 ;
        RECT 372.720 792.960 374.640 793.365 ;
        RECT 375.480 792.960 377.860 793.365 ;
        RECT 378.700 792.960 381.080 793.365 ;
        RECT 381.920 792.960 384.300 793.365 ;
        RECT 385.140 792.960 387.060 793.365 ;
        RECT 387.900 792.960 390.280 793.365 ;
        RECT 391.120 792.960 393.500 793.365 ;
        RECT 394.340 792.960 396.260 793.365 ;
        RECT 397.100 792.960 399.480 793.365 ;
        RECT 400.320 792.960 402.700 793.365 ;
        RECT 403.540 792.960 405.460 793.365 ;
        RECT 406.300 792.960 408.680 793.365 ;
        RECT 409.520 792.960 411.900 793.365 ;
        RECT 412.740 792.960 414.660 793.365 ;
        RECT 415.500 792.960 417.880 793.365 ;
        RECT 418.720 792.960 421.100 793.365 ;
        RECT 421.940 792.960 424.320 793.365 ;
        RECT 425.160 792.960 427.080 793.365 ;
        RECT 427.920 792.960 430.300 793.365 ;
        RECT 431.140 792.960 433.520 793.365 ;
        RECT 434.360 792.960 436.280 793.365 ;
        RECT 437.120 792.960 439.500 793.365 ;
        RECT 440.340 792.960 442.720 793.365 ;
        RECT 443.560 792.960 445.480 793.365 ;
        RECT 446.320 792.960 448.700 793.365 ;
        RECT 449.540 792.960 451.920 793.365 ;
        RECT 452.760 792.960 454.680 793.365 ;
        RECT 455.520 792.960 457.900 793.365 ;
        RECT 458.740 792.960 461.120 793.365 ;
        RECT 461.960 792.960 463.880 793.365 ;
        RECT 464.720 792.960 467.100 793.365 ;
        RECT 467.940 792.960 470.320 793.365 ;
        RECT 471.160 792.960 473.540 793.365 ;
        RECT 474.380 792.960 476.300 793.365 ;
        RECT 477.140 792.960 479.520 793.365 ;
        RECT 480.360 792.960 482.740 793.365 ;
        RECT 483.580 792.960 485.500 793.365 ;
        RECT 486.340 792.960 488.720 793.365 ;
        RECT 489.560 792.960 491.940 793.365 ;
        RECT 492.780 792.960 494.700 793.365 ;
        RECT 495.540 792.960 497.920 793.365 ;
        RECT 498.760 792.960 501.140 793.365 ;
        RECT 501.980 792.960 503.900 793.365 ;
        RECT 504.740 792.960 507.120 793.365 ;
        RECT 507.960 792.960 510.340 793.365 ;
        RECT 511.180 792.960 513.100 793.365 ;
        RECT 513.940 792.960 516.320 793.365 ;
        RECT 517.160 792.960 519.540 793.365 ;
        RECT 520.380 792.960 522.760 793.365 ;
        RECT 523.600 792.960 525.520 793.365 ;
        RECT 526.360 792.960 528.740 793.365 ;
        RECT 529.580 792.960 531.960 793.365 ;
        RECT 532.800 792.960 534.720 793.365 ;
        RECT 535.560 792.960 537.940 793.365 ;
        RECT 538.780 792.960 541.160 793.365 ;
        RECT 542.000 792.960 543.920 793.365 ;
        RECT 544.760 792.960 547.140 793.365 ;
        RECT 547.980 792.960 550.360 793.365 ;
        RECT 551.200 792.960 553.120 793.365 ;
        RECT 553.960 792.960 556.340 793.365 ;
        RECT 557.180 792.960 559.560 793.365 ;
        RECT 560.400 792.960 562.320 793.365 ;
        RECT 563.160 792.960 565.540 793.365 ;
        RECT 566.380 792.960 568.760 793.365 ;
        RECT 569.600 792.960 571.980 793.365 ;
        RECT 572.820 792.960 574.740 793.365 ;
        RECT 575.580 792.960 577.960 793.365 ;
        RECT 578.800 792.960 581.180 793.365 ;
        RECT 582.020 792.960 583.940 793.365 ;
        RECT 584.780 792.960 587.160 793.365 ;
        RECT 588.000 792.960 590.380 793.365 ;
        RECT 591.220 792.960 593.140 793.365 ;
        RECT 593.980 792.960 596.360 793.365 ;
        RECT 597.200 792.960 599.580 793.365 ;
        RECT 600.420 792.960 602.340 793.365 ;
        RECT 603.180 792.960 605.560 793.365 ;
        RECT 606.400 792.960 608.780 793.365 ;
        RECT 609.620 792.960 612.000 793.365 ;
        RECT 612.840 792.960 614.760 793.365 ;
        RECT 615.600 792.960 617.980 793.365 ;
        RECT 618.820 792.960 621.200 793.365 ;
        RECT 622.040 792.960 623.960 793.365 ;
        RECT 624.800 792.960 627.180 793.365 ;
        RECT 628.020 792.960 630.400 793.365 ;
        RECT 631.240 792.960 633.160 793.365 ;
        RECT 634.000 792.960 636.380 793.365 ;
        RECT 637.220 792.960 639.600 793.365 ;
        RECT 640.440 792.960 642.360 793.365 ;
        RECT 643.200 792.960 645.580 793.365 ;
        RECT 646.420 792.960 648.800 793.365 ;
        RECT 649.640 792.960 651.560 793.365 ;
        RECT 652.400 792.960 654.780 793.365 ;
        RECT 655.620 792.960 658.000 793.365 ;
        RECT 658.840 792.960 661.220 793.365 ;
        RECT 662.060 792.960 663.980 793.365 ;
        RECT 664.820 792.960 667.200 793.365 ;
        RECT 668.040 792.960 670.420 793.365 ;
        RECT 671.260 792.960 673.180 793.365 ;
        RECT 674.020 792.960 676.400 793.365 ;
        RECT 677.240 792.960 679.620 793.365 ;
        RECT 680.460 792.960 682.380 793.365 ;
        RECT 683.220 792.960 685.600 793.365 ;
        RECT 686.440 792.960 688.820 793.365 ;
        RECT 689.660 792.960 691.580 793.365 ;
        RECT 692.420 792.960 694.800 793.365 ;
        RECT 695.640 792.960 698.020 793.365 ;
        RECT 698.860 792.960 700.780 793.365 ;
        RECT 701.620 792.960 704.000 793.365 ;
        RECT 704.840 792.960 707.220 793.365 ;
        RECT 708.060 792.960 710.440 793.365 ;
        RECT 711.280 792.960 713.200 793.365 ;
        RECT 714.040 792.960 716.420 793.365 ;
        RECT 717.260 792.960 719.640 793.365 ;
        RECT 720.480 792.960 722.400 793.365 ;
        RECT 723.240 792.960 725.620 793.365 ;
        RECT 726.460 792.960 728.840 793.365 ;
        RECT 729.680 792.960 731.600 793.365 ;
        RECT 732.440 792.960 734.820 793.365 ;
        RECT 735.660 792.960 738.040 793.365 ;
        RECT 738.880 792.960 740.800 793.365 ;
        RECT 741.640 792.960 744.020 793.365 ;
        RECT 744.860 792.960 747.240 793.365 ;
        RECT 748.080 792.960 750.000 793.365 ;
        RECT 750.840 792.960 753.220 793.365 ;
        RECT 754.060 792.960 756.440 793.365 ;
        RECT 757.280 792.960 759.660 793.365 ;
        RECT 760.500 792.960 762.420 793.365 ;
        RECT 763.260 792.960 765.640 793.365 ;
        RECT 766.480 792.960 768.860 793.365 ;
        RECT 769.700 792.960 771.620 793.365 ;
        RECT 772.460 792.960 774.840 793.365 ;
        RECT 775.680 792.960 778.060 793.365 ;
        RECT 778.900 792.960 780.820 793.365 ;
        RECT 781.660 792.960 784.040 793.365 ;
        RECT 784.880 792.960 787.260 793.365 ;
        RECT 788.100 792.960 790.020 793.365 ;
        RECT 790.860 792.960 793.240 793.365 ;
        RECT 794.080 792.960 796.460 793.365 ;
        RECT 0.030 0.115 797.010 792.960 ;
      LAYER met3 ;
        RECT 6.895 792.480 794.150 793.345 ;
        RECT 6.895 787.760 795.205 792.480 ;
        RECT 6.895 786.360 794.150 787.760 ;
        RECT 6.895 781.640 795.205 786.360 ;
        RECT 6.895 780.240 794.150 781.640 ;
        RECT 6.895 775.520 795.205 780.240 ;
        RECT 6.895 774.120 794.150 775.520 ;
        RECT 6.895 769.400 795.205 774.120 ;
        RECT 6.895 768.000 794.150 769.400 ;
        RECT 6.895 763.280 795.205 768.000 ;
        RECT 6.895 761.880 794.150 763.280 ;
        RECT 6.895 757.160 795.205 761.880 ;
        RECT 6.895 755.760 794.150 757.160 ;
        RECT 6.895 751.040 795.205 755.760 ;
        RECT 6.895 749.640 794.150 751.040 ;
        RECT 6.895 744.920 795.205 749.640 ;
        RECT 6.895 743.520 794.150 744.920 ;
        RECT 6.895 738.800 795.205 743.520 ;
        RECT 6.895 737.400 794.150 738.800 ;
        RECT 6.895 732.680 795.205 737.400 ;
        RECT 6.895 731.280 794.150 732.680 ;
        RECT 6.895 726.560 795.205 731.280 ;
        RECT 6.895 725.160 794.150 726.560 ;
        RECT 6.895 720.440 795.205 725.160 ;
        RECT 6.895 719.040 794.150 720.440 ;
        RECT 6.895 714.320 795.205 719.040 ;
        RECT 6.895 712.920 794.150 714.320 ;
        RECT 6.895 708.200 795.205 712.920 ;
        RECT 6.895 706.800 794.150 708.200 ;
        RECT 6.895 702.080 795.205 706.800 ;
        RECT 6.895 700.680 794.150 702.080 ;
        RECT 6.895 695.960 795.205 700.680 ;
        RECT 6.895 694.560 794.150 695.960 ;
        RECT 6.895 689.840 795.205 694.560 ;
        RECT 6.895 688.440 794.150 689.840 ;
        RECT 6.895 683.720 795.205 688.440 ;
        RECT 6.895 682.320 794.150 683.720 ;
        RECT 6.895 677.600 795.205 682.320 ;
        RECT 6.895 676.200 794.150 677.600 ;
        RECT 6.895 671.480 795.205 676.200 ;
        RECT 6.895 670.080 794.150 671.480 ;
        RECT 6.895 664.680 795.205 670.080 ;
        RECT 6.895 663.280 794.150 664.680 ;
        RECT 6.895 658.560 795.205 663.280 ;
        RECT 6.895 657.160 794.150 658.560 ;
        RECT 6.895 652.440 795.205 657.160 ;
        RECT 6.895 651.040 794.150 652.440 ;
        RECT 6.895 646.320 795.205 651.040 ;
        RECT 6.895 644.920 794.150 646.320 ;
        RECT 6.895 640.200 795.205 644.920 ;
        RECT 6.895 638.800 794.150 640.200 ;
        RECT 6.895 634.080 795.205 638.800 ;
        RECT 6.895 632.680 794.150 634.080 ;
        RECT 6.895 627.960 795.205 632.680 ;
        RECT 6.895 626.560 794.150 627.960 ;
        RECT 6.895 621.840 795.205 626.560 ;
        RECT 6.895 620.440 794.150 621.840 ;
        RECT 6.895 615.720 795.205 620.440 ;
        RECT 6.895 614.320 794.150 615.720 ;
        RECT 6.895 609.600 795.205 614.320 ;
        RECT 6.895 608.200 794.150 609.600 ;
        RECT 6.895 603.480 795.205 608.200 ;
        RECT 6.895 602.080 794.150 603.480 ;
        RECT 6.895 597.360 795.205 602.080 ;
        RECT 6.895 595.960 794.150 597.360 ;
        RECT 6.895 591.240 795.205 595.960 ;
        RECT 6.895 589.840 794.150 591.240 ;
        RECT 6.895 585.120 795.205 589.840 ;
        RECT 6.895 583.720 794.150 585.120 ;
        RECT 6.895 579.000 795.205 583.720 ;
        RECT 6.895 577.600 794.150 579.000 ;
        RECT 6.895 572.880 795.205 577.600 ;
        RECT 6.895 571.480 794.150 572.880 ;
        RECT 6.895 566.760 795.205 571.480 ;
        RECT 6.895 565.360 794.150 566.760 ;
        RECT 6.895 560.640 795.205 565.360 ;
        RECT 6.895 559.240 794.150 560.640 ;
        RECT 6.895 554.520 795.205 559.240 ;
        RECT 6.895 553.120 794.150 554.520 ;
        RECT 6.895 548.400 795.205 553.120 ;
        RECT 6.895 547.000 794.150 548.400 ;
        RECT 6.895 542.280 795.205 547.000 ;
        RECT 6.895 540.880 794.150 542.280 ;
        RECT 6.895 536.160 795.205 540.880 ;
        RECT 6.895 534.760 794.150 536.160 ;
        RECT 6.895 529.360 795.205 534.760 ;
        RECT 6.895 527.960 794.150 529.360 ;
        RECT 6.895 523.240 795.205 527.960 ;
        RECT 6.895 521.840 794.150 523.240 ;
        RECT 6.895 517.120 795.205 521.840 ;
        RECT 6.895 515.720 794.150 517.120 ;
        RECT 6.895 511.000 795.205 515.720 ;
        RECT 6.895 509.600 794.150 511.000 ;
        RECT 6.895 504.880 795.205 509.600 ;
        RECT 6.895 503.480 794.150 504.880 ;
        RECT 6.895 498.760 795.205 503.480 ;
        RECT 6.895 497.360 794.150 498.760 ;
        RECT 6.895 492.640 795.205 497.360 ;
        RECT 6.895 491.240 794.150 492.640 ;
        RECT 6.895 486.520 795.205 491.240 ;
        RECT 6.895 485.120 794.150 486.520 ;
        RECT 6.895 480.400 795.205 485.120 ;
        RECT 6.895 479.000 794.150 480.400 ;
        RECT 6.895 474.280 795.205 479.000 ;
        RECT 6.895 472.880 794.150 474.280 ;
        RECT 6.895 468.160 795.205 472.880 ;
        RECT 6.895 466.760 794.150 468.160 ;
        RECT 6.895 462.040 795.205 466.760 ;
        RECT 6.895 460.640 794.150 462.040 ;
        RECT 6.895 455.920 795.205 460.640 ;
        RECT 6.895 454.520 794.150 455.920 ;
        RECT 6.895 449.800 795.205 454.520 ;
        RECT 6.895 448.400 794.150 449.800 ;
        RECT 6.895 443.680 795.205 448.400 ;
        RECT 6.895 442.280 794.150 443.680 ;
        RECT 6.895 437.560 795.205 442.280 ;
        RECT 6.895 436.160 794.150 437.560 ;
        RECT 6.895 431.440 795.205 436.160 ;
        RECT 6.895 430.040 794.150 431.440 ;
        RECT 6.895 425.320 795.205 430.040 ;
        RECT 6.895 423.920 794.150 425.320 ;
        RECT 6.895 419.200 795.205 423.920 ;
        RECT 6.895 417.800 794.150 419.200 ;
        RECT 6.895 413.080 795.205 417.800 ;
        RECT 6.895 411.680 794.150 413.080 ;
        RECT 6.895 406.960 795.205 411.680 ;
        RECT 6.895 405.560 794.150 406.960 ;
        RECT 6.895 400.840 795.205 405.560 ;
        RECT 6.895 399.440 794.150 400.840 ;
        RECT 6.895 394.040 795.205 399.440 ;
        RECT 6.895 392.640 794.150 394.040 ;
        RECT 6.895 387.920 795.205 392.640 ;
        RECT 6.895 386.520 794.150 387.920 ;
        RECT 6.895 381.800 795.205 386.520 ;
        RECT 6.895 380.400 794.150 381.800 ;
        RECT 6.895 375.680 795.205 380.400 ;
        RECT 6.895 374.280 794.150 375.680 ;
        RECT 6.895 369.560 795.205 374.280 ;
        RECT 6.895 368.160 794.150 369.560 ;
        RECT 6.895 363.440 795.205 368.160 ;
        RECT 6.895 362.040 794.150 363.440 ;
        RECT 6.895 357.320 795.205 362.040 ;
        RECT 6.895 355.920 794.150 357.320 ;
        RECT 6.895 351.200 795.205 355.920 ;
        RECT 6.895 349.800 794.150 351.200 ;
        RECT 6.895 345.080 795.205 349.800 ;
        RECT 6.895 343.680 794.150 345.080 ;
        RECT 6.895 338.960 795.205 343.680 ;
        RECT 6.895 337.560 794.150 338.960 ;
        RECT 6.895 332.840 795.205 337.560 ;
        RECT 6.895 331.440 794.150 332.840 ;
        RECT 6.895 326.720 795.205 331.440 ;
        RECT 6.895 325.320 794.150 326.720 ;
        RECT 6.895 320.600 795.205 325.320 ;
        RECT 6.895 319.200 794.150 320.600 ;
        RECT 6.895 314.480 795.205 319.200 ;
        RECT 6.895 313.080 794.150 314.480 ;
        RECT 6.895 308.360 795.205 313.080 ;
        RECT 6.895 306.960 794.150 308.360 ;
        RECT 6.895 302.240 795.205 306.960 ;
        RECT 6.895 300.840 794.150 302.240 ;
        RECT 6.895 296.120 795.205 300.840 ;
        RECT 6.895 294.720 794.150 296.120 ;
        RECT 6.895 290.000 795.205 294.720 ;
        RECT 6.895 288.600 794.150 290.000 ;
        RECT 6.895 283.880 795.205 288.600 ;
        RECT 6.895 282.480 794.150 283.880 ;
        RECT 6.895 277.760 795.205 282.480 ;
        RECT 6.895 276.360 794.150 277.760 ;
        RECT 6.895 271.640 795.205 276.360 ;
        RECT 6.895 270.240 794.150 271.640 ;
        RECT 6.895 264.840 795.205 270.240 ;
        RECT 6.895 263.440 794.150 264.840 ;
        RECT 6.895 258.720 795.205 263.440 ;
        RECT 6.895 257.320 794.150 258.720 ;
        RECT 6.895 252.600 795.205 257.320 ;
        RECT 6.895 251.200 794.150 252.600 ;
        RECT 6.895 246.480 795.205 251.200 ;
        RECT 6.895 245.080 794.150 246.480 ;
        RECT 6.895 240.360 795.205 245.080 ;
        RECT 6.895 238.960 794.150 240.360 ;
        RECT 6.895 234.240 795.205 238.960 ;
        RECT 6.895 232.840 794.150 234.240 ;
        RECT 6.895 228.120 795.205 232.840 ;
        RECT 6.895 226.720 794.150 228.120 ;
        RECT 6.895 222.000 795.205 226.720 ;
        RECT 6.895 220.600 794.150 222.000 ;
        RECT 6.895 215.880 795.205 220.600 ;
        RECT 6.895 214.480 794.150 215.880 ;
        RECT 6.895 209.760 795.205 214.480 ;
        RECT 6.895 208.360 794.150 209.760 ;
        RECT 6.895 203.640 795.205 208.360 ;
        RECT 6.895 202.240 794.150 203.640 ;
        RECT 6.895 197.520 795.205 202.240 ;
        RECT 6.895 196.120 794.150 197.520 ;
        RECT 6.895 191.400 795.205 196.120 ;
        RECT 6.895 190.000 794.150 191.400 ;
        RECT 6.895 185.280 795.205 190.000 ;
        RECT 6.895 183.880 794.150 185.280 ;
        RECT 6.895 179.160 795.205 183.880 ;
        RECT 6.895 177.760 794.150 179.160 ;
        RECT 6.895 173.040 795.205 177.760 ;
        RECT 6.895 171.640 794.150 173.040 ;
        RECT 6.895 166.920 795.205 171.640 ;
        RECT 6.895 165.520 794.150 166.920 ;
        RECT 6.895 160.800 795.205 165.520 ;
        RECT 6.895 159.400 794.150 160.800 ;
        RECT 6.895 154.680 795.205 159.400 ;
        RECT 6.895 153.280 794.150 154.680 ;
        RECT 6.895 148.560 795.205 153.280 ;
        RECT 6.895 147.160 794.150 148.560 ;
        RECT 6.895 142.440 795.205 147.160 ;
        RECT 6.895 141.040 794.150 142.440 ;
        RECT 6.895 136.320 795.205 141.040 ;
        RECT 6.895 134.920 794.150 136.320 ;
        RECT 6.895 129.520 795.205 134.920 ;
        RECT 6.895 128.120 794.150 129.520 ;
        RECT 6.895 123.400 795.205 128.120 ;
        RECT 6.895 122.000 794.150 123.400 ;
        RECT 6.895 117.280 795.205 122.000 ;
        RECT 6.895 115.880 794.150 117.280 ;
        RECT 6.895 111.160 795.205 115.880 ;
        RECT 6.895 109.760 794.150 111.160 ;
        RECT 6.895 105.040 795.205 109.760 ;
        RECT 6.895 103.640 794.150 105.040 ;
        RECT 6.895 98.920 795.205 103.640 ;
        RECT 6.895 97.520 794.150 98.920 ;
        RECT 6.895 92.800 795.205 97.520 ;
        RECT 6.895 91.400 794.150 92.800 ;
        RECT 6.895 86.680 795.205 91.400 ;
        RECT 6.895 85.280 794.150 86.680 ;
        RECT 6.895 80.560 795.205 85.280 ;
        RECT 6.895 79.160 794.150 80.560 ;
        RECT 6.895 74.440 795.205 79.160 ;
        RECT 6.895 73.040 794.150 74.440 ;
        RECT 6.895 68.320 795.205 73.040 ;
        RECT 6.895 66.920 794.150 68.320 ;
        RECT 6.895 62.200 795.205 66.920 ;
        RECT 6.895 60.800 794.150 62.200 ;
        RECT 6.895 56.080 795.205 60.800 ;
        RECT 6.895 54.680 794.150 56.080 ;
        RECT 6.895 49.960 795.205 54.680 ;
        RECT 6.895 48.560 794.150 49.960 ;
        RECT 6.895 43.840 795.205 48.560 ;
        RECT 6.895 42.440 794.150 43.840 ;
        RECT 6.895 37.720 795.205 42.440 ;
        RECT 6.895 36.320 794.150 37.720 ;
        RECT 6.895 31.600 795.205 36.320 ;
        RECT 6.895 30.200 794.150 31.600 ;
        RECT 6.895 25.480 795.205 30.200 ;
        RECT 6.895 24.080 794.150 25.480 ;
        RECT 6.895 19.360 795.205 24.080 ;
        RECT 6.895 17.960 794.150 19.360 ;
        RECT 6.895 13.240 795.205 17.960 ;
        RECT 6.895 11.840 794.150 13.240 ;
        RECT 6.895 7.120 795.205 11.840 ;
        RECT 6.895 5.720 794.150 7.120 ;
        RECT 6.895 1.000 795.205 5.720 ;
        RECT 6.895 0.135 794.150 1.000 ;
      LAYER met4 ;
        RECT 14.485 20.535 19.190 786.545 ;
        RECT 21.590 786.440 95.990 786.545 ;
        RECT 21.590 20.535 22.490 786.440 ;
        RECT 24.890 20.535 25.790 786.440 ;
        RECT 28.190 20.535 29.090 786.440 ;
        RECT 31.490 20.535 95.990 786.440 ;
        RECT 98.390 786.440 172.790 786.545 ;
        RECT 98.390 20.535 99.290 786.440 ;
        RECT 101.690 20.535 102.590 786.440 ;
        RECT 104.990 20.535 105.890 786.440 ;
        RECT 108.290 20.535 172.790 786.440 ;
        RECT 175.190 786.440 249.590 786.545 ;
        RECT 175.190 20.535 176.090 786.440 ;
        RECT 178.490 20.535 179.390 786.440 ;
        RECT 181.790 20.535 182.690 786.440 ;
        RECT 185.090 20.535 249.590 786.440 ;
        RECT 251.990 786.440 326.390 786.545 ;
        RECT 251.990 20.535 252.890 786.440 ;
        RECT 255.290 20.535 256.190 786.440 ;
        RECT 258.590 20.535 259.490 786.440 ;
        RECT 261.890 20.535 326.390 786.440 ;
        RECT 328.790 786.440 403.190 786.545 ;
        RECT 328.790 20.535 329.690 786.440 ;
        RECT 332.090 20.535 332.990 786.440 ;
        RECT 335.390 20.535 336.290 786.440 ;
        RECT 338.690 20.535 403.190 786.440 ;
        RECT 405.590 786.440 479.990 786.545 ;
        RECT 405.590 20.535 406.490 786.440 ;
        RECT 408.890 20.535 409.790 786.440 ;
        RECT 412.190 20.535 413.090 786.440 ;
        RECT 415.490 20.535 479.990 786.440 ;
        RECT 482.390 786.440 556.790 786.545 ;
        RECT 482.390 20.535 483.290 786.440 ;
        RECT 485.690 20.535 486.590 786.440 ;
        RECT 488.990 20.535 489.890 786.440 ;
        RECT 492.290 20.535 556.790 786.440 ;
        RECT 559.190 786.440 633.590 786.545 ;
        RECT 559.190 20.535 560.090 786.440 ;
        RECT 562.490 20.535 563.390 786.440 ;
        RECT 565.790 20.535 566.690 786.440 ;
        RECT 569.090 20.535 633.590 786.440 ;
        RECT 635.990 786.440 710.390 786.545 ;
        RECT 635.990 20.535 636.890 786.440 ;
        RECT 639.290 20.535 640.190 786.440 ;
        RECT 642.590 20.535 643.490 786.440 ;
        RECT 645.890 20.535 710.390 786.440 ;
        RECT 712.790 786.440 786.695 786.545 ;
        RECT 712.790 20.535 713.690 786.440 ;
        RECT 716.090 20.535 716.990 786.440 ;
        RECT 719.390 20.535 720.290 786.440 ;
        RECT 722.690 20.535 786.695 786.440 ;
  END
END multiply_4
END LIBRARY

