VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dcache
  CLASS BLOCK ;
  FOREIGN dcache ;
  ORIGIN 0.000 0.000 ;
  SIZE 717.990 BY 720.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END clk
  PIN d_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END d_in[0]
  PIN d_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END d_in[100]
  PIN d_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END d_in[101]
  PIN d_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END d_in[102]
  PIN d_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END d_in[103]
  PIN d_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 4.000 ;
    END
  END d_in[104]
  PIN d_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 0.000 361.470 4.000 ;
    END
  END d_in[105]
  PIN d_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END d_in[106]
  PIN d_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END d_in[107]
  PIN d_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END d_in[108]
  PIN d_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END d_in[109]
  PIN d_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END d_in[10]
  PIN d_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END d_in[110]
  PIN d_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 0.000 381.710 4.000 ;
    END
  END d_in[111]
  PIN d_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END d_in[112]
  PIN d_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END d_in[113]
  PIN d_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 0.000 391.830 4.000 ;
    END
  END d_in[114]
  PIN d_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 0.000 395.510 4.000 ;
    END
  END d_in[115]
  PIN d_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END d_in[116]
  PIN d_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 0.000 402.410 4.000 ;
    END
  END d_in[117]
  PIN d_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.350 0.000 405.630 4.000 ;
    END
  END d_in[118]
  PIN d_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END d_in[119]
  PIN d_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END d_in[11]
  PIN d_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END d_in[120]
  PIN d_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END d_in[121]
  PIN d_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END d_in[122]
  PIN d_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 0.000 422.650 4.000 ;
    END
  END d_in[123]
  PIN d_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 0.000 425.870 4.000 ;
    END
  END d_in[124]
  PIN d_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 0.000 429.550 4.000 ;
    END
  END d_in[125]
  PIN d_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END d_in[126]
  PIN d_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 0.000 435.990 4.000 ;
    END
  END d_in[127]
  PIN d_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 0.000 439.670 4.000 ;
    END
  END d_in[128]
  PIN d_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 0.000 442.890 4.000 ;
    END
  END d_in[129]
  PIN d_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END d_in[12]
  PIN d_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 4.000 ;
    END
  END d_in[130]
  PIN d_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END d_in[131]
  PIN d_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 0.000 453.010 4.000 ;
    END
  END d_in[132]
  PIN d_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 4.000 ;
    END
  END d_in[133]
  PIN d_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.630 0.000 459.910 4.000 ;
    END
  END d_in[134]
  PIN d_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 0.000 463.130 4.000 ;
    END
  END d_in[135]
  PIN d_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 0.000 466.810 4.000 ;
    END
  END d_in[136]
  PIN d_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 0.000 470.030 4.000 ;
    END
  END d_in[137]
  PIN d_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END d_in[138]
  PIN d_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END d_in[139]
  PIN d_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END d_in[13]
  PIN d_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END d_in[140]
  PIN d_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 0.000 483.830 4.000 ;
    END
  END d_in[141]
  PIN d_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 0.000 487.050 4.000 ;
    END
  END d_in[142]
  PIN d_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 4.000 ;
    END
  END d_in[14]
  PIN d_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END d_in[15]
  PIN d_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END d_in[16]
  PIN d_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END d_in[17]
  PIN d_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END d_in[18]
  PIN d_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END d_in[19]
  PIN d_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END d_in[1]
  PIN d_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END d_in[20]
  PIN d_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END d_in[21]
  PIN d_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END d_in[22]
  PIN d_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END d_in[23]
  PIN d_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END d_in[24]
  PIN d_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END d_in[25]
  PIN d_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END d_in[26]
  PIN d_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END d_in[27]
  PIN d_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END d_in[28]
  PIN d_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END d_in[29]
  PIN d_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END d_in[2]
  PIN d_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END d_in[30]
  PIN d_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END d_in[31]
  PIN d_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END d_in[32]
  PIN d_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END d_in[33]
  PIN d_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END d_in[34]
  PIN d_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END d_in[35]
  PIN d_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END d_in[36]
  PIN d_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END d_in[37]
  PIN d_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END d_in[38]
  PIN d_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END d_in[39]
  PIN d_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END d_in[3]
  PIN d_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END d_in[40]
  PIN d_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END d_in[41]
  PIN d_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END d_in[42]
  PIN d_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END d_in[43]
  PIN d_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END d_in[44]
  PIN d_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END d_in[45]
  PIN d_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END d_in[46]
  PIN d_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END d_in[47]
  PIN d_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END d_in[48]
  PIN d_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END d_in[49]
  PIN d_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END d_in[4]
  PIN d_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END d_in[50]
  PIN d_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END d_in[51]
  PIN d_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END d_in[52]
  PIN d_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 4.000 ;
    END
  END d_in[53]
  PIN d_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END d_in[54]
  PIN d_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END d_in[55]
  PIN d_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 4.000 ;
    END
  END d_in[56]
  PIN d_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END d_in[57]
  PIN d_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END d_in[58]
  PIN d_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 0.000 205.070 4.000 ;
    END
  END d_in[59]
  PIN d_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 4.000 ;
    END
  END d_in[5]
  PIN d_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END d_in[60]
  PIN d_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END d_in[61]
  PIN d_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END d_in[62]
  PIN d_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END d_in[63]
  PIN d_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END d_in[64]
  PIN d_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END d_in[65]
  PIN d_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END d_in[66]
  PIN d_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END d_in[67]
  PIN d_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END d_in[68]
  PIN d_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 0.000 239.110 4.000 ;
    END
  END d_in[69]
  PIN d_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END d_in[6]
  PIN d_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 4.000 ;
    END
  END d_in[70]
  PIN d_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END d_in[71]
  PIN d_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END d_in[72]
  PIN d_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 0.000 252.910 4.000 ;
    END
  END d_in[73]
  PIN d_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END d_in[74]
  PIN d_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END d_in[75]
  PIN d_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END d_in[76]
  PIN d_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 0.000 266.250 4.000 ;
    END
  END d_in[77]
  PIN d_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END d_in[78]
  PIN d_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END d_in[79]
  PIN d_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END d_in[7]
  PIN d_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END d_in[80]
  PIN d_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END d_in[81]
  PIN d_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 4.000 ;
    END
  END d_in[82]
  PIN d_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END d_in[83]
  PIN d_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END d_in[84]
  PIN d_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END d_in[85]
  PIN d_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END d_in[86]
  PIN d_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 4.000 ;
    END
  END d_in[87]
  PIN d_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END d_in[88]
  PIN d_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END d_in[89]
  PIN d_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END d_in[8]
  PIN d_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 0.000 310.410 4.000 ;
    END
  END d_in[90]
  PIN d_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END d_in[91]
  PIN d_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 0.000 317.310 4.000 ;
    END
  END d_in[92]
  PIN d_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 4.000 ;
    END
  END d_in[93]
  PIN d_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END d_in[94]
  PIN d_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END d_in[95]
  PIN d_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 4.000 ;
    END
  END d_in[96]
  PIN d_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END d_in[97]
  PIN d_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END d_in[98]
  PIN d_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 4.000 ;
    END
  END d_in[99]
  PIN d_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END d_in[9]
  PIN d_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.450 0.000 490.730 4.000 ;
    END
  END d_out[0]
  PIN d_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 0.000 524.310 4.000 ;
    END
  END d_out[10]
  PIN d_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 0.000 527.990 4.000 ;
    END
  END d_out[11]
  PIN d_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.930 0.000 531.210 4.000 ;
    END
  END d_out[12]
  PIN d_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 0.000 534.430 4.000 ;
    END
  END d_out[13]
  PIN d_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END d_out[14]
  PIN d_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END d_out[15]
  PIN d_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 0.000 545.010 4.000 ;
    END
  END d_out[16]
  PIN d_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 0.000 548.230 4.000 ;
    END
  END d_out[17]
  PIN d_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 0.000 551.450 4.000 ;
    END
  END d_out[18]
  PIN d_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.850 0.000 555.130 4.000 ;
    END
  END d_out[19]
  PIN d_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.670 0.000 493.950 4.000 ;
    END
  END d_out[1]
  PIN d_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.070 0.000 558.350 4.000 ;
    END
  END d_out[20]
  PIN d_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 0.000 562.030 4.000 ;
    END
  END d_out[21]
  PIN d_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 0.000 565.250 4.000 ;
    END
  END d_out[22]
  PIN d_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.190 0.000 568.470 4.000 ;
    END
  END d_out[23]
  PIN d_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.870 0.000 572.150 4.000 ;
    END
  END d_out[24]
  PIN d_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.090 0.000 575.370 4.000 ;
    END
  END d_out[25]
  PIN d_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 0.000 578.590 4.000 ;
    END
  END d_out[26]
  PIN d_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 0.000 582.270 4.000 ;
    END
  END d_out[27]
  PIN d_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END d_out[28]
  PIN d_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 0.000 589.170 4.000 ;
    END
  END d_out[29]
  PIN d_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END d_out[2]
  PIN d_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 0.000 592.390 4.000 ;
    END
  END d_out[30]
  PIN d_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 4.000 ;
    END
  END d_out[31]
  PIN d_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END d_out[32]
  PIN d_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 0.000 602.510 4.000 ;
    END
  END d_out[33]
  PIN d_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 0.000 606.190 4.000 ;
    END
  END d_out[34]
  PIN d_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 0.000 609.410 4.000 ;
    END
  END d_out[35]
  PIN d_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 0.000 612.630 4.000 ;
    END
  END d_out[36]
  PIN d_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.030 0.000 616.310 4.000 ;
    END
  END d_out[37]
  PIN d_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.250 0.000 619.530 4.000 ;
    END
  END d_out[38]
  PIN d_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 0.000 622.750 4.000 ;
    END
  END d_out[39]
  PIN d_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 0.000 500.850 4.000 ;
    END
  END d_out[3]
  PIN d_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.150 0.000 626.430 4.000 ;
    END
  END d_out[40]
  PIN d_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.370 0.000 629.650 4.000 ;
    END
  END d_out[41]
  PIN d_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.050 0.000 633.330 4.000 ;
    END
  END d_out[42]
  PIN d_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 0.000 636.550 4.000 ;
    END
  END d_out[43]
  PIN d_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.490 0.000 639.770 4.000 ;
    END
  END d_out[44]
  PIN d_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 0.000 643.450 4.000 ;
    END
  END d_out[45]
  PIN d_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 0.000 646.670 4.000 ;
    END
  END d_out[46]
  PIN d_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 0.000 649.890 4.000 ;
    END
  END d_out[47]
  PIN d_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 4.000 ;
    END
  END d_out[48]
  PIN d_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 0.000 656.790 4.000 ;
    END
  END d_out[49]
  PIN d_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 0.000 504.070 4.000 ;
    END
  END d_out[4]
  PIN d_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END d_out[50]
  PIN d_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END d_out[51]
  PIN d_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END d_out[52]
  PIN d_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 0.000 670.590 4.000 ;
    END
  END d_out[53]
  PIN d_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 0.000 673.810 4.000 ;
    END
  END d_out[54]
  PIN d_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.210 0.000 677.490 4.000 ;
    END
  END d_out[55]
  PIN d_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 0.000 680.710 4.000 ;
    END
  END d_out[56]
  PIN d_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.650 0.000 683.930 4.000 ;
    END
  END d_out[57]
  PIN d_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.330 0.000 687.610 4.000 ;
    END
  END d_out[58]
  PIN d_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.550 0.000 690.830 4.000 ;
    END
  END d_out[59]
  PIN d_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.010 0.000 507.290 4.000 ;
    END
  END d_out[5]
  PIN d_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 0.000 694.050 4.000 ;
    END
  END d_out[60]
  PIN d_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 0.000 697.730 4.000 ;
    END
  END d_out[61]
  PIN d_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.670 0.000 700.950 4.000 ;
    END
  END d_out[62]
  PIN d_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.350 0.000 704.630 4.000 ;
    END
  END d_out[63]
  PIN d_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 0.000 707.850 4.000 ;
    END
  END d_out[64]
  PIN d_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.790 0.000 711.070 4.000 ;
    END
  END d_out[65]
  PIN d_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.470 0.000 714.750 4.000 ;
    END
  END d_out[66]
  PIN d_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 0.000 717.970 4.000 ;
    END
  END d_out[67]
  PIN d_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 0.000 510.970 4.000 ;
    END
  END d_out[6]
  PIN d_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 0.000 514.190 4.000 ;
    END
  END d_out[7]
  PIN d_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 0.000 517.870 4.000 ;
    END
  END d_out[8]
  PIN d_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 0.000 521.090 4.000 ;
    END
  END d_out[9]
  PIN m_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END m_in[0]
  PIN m_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.560 4.000 367.160 ;
    END
  END m_in[100]
  PIN m_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END m_in[101]
  PIN m_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 373.360 4.000 373.960 ;
    END
  END m_in[102]
  PIN m_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END m_in[103]
  PIN m_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END m_in[104]
  PIN m_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END m_in[105]
  PIN m_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 388.320 4.000 388.920 ;
    END
  END m_in[106]
  PIN m_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END m_in[107]
  PIN m_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.120 4.000 395.720 ;
    END
  END m_in[108]
  PIN m_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END m_in[109]
  PIN m_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END m_in[10]
  PIN m_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END m_in[110]
  PIN m_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.000 4.000 406.600 ;
    END
  END m_in[111]
  PIN m_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END m_in[112]
  PIN m_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.800 4.000 413.400 ;
    END
  END m_in[113]
  PIN m_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.880 4.000 417.480 ;
    END
  END m_in[114]
  PIN m_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END m_in[115]
  PIN m_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.680 4.000 424.280 ;
    END
  END m_in[116]
  PIN m_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END m_in[117]
  PIN m_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END m_in[118]
  PIN m_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 434.560 4.000 435.160 ;
    END
  END m_in[119]
  PIN m_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END m_in[11]
  PIN m_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END m_in[120]
  PIN m_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END m_in[121]
  PIN m_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END m_in[122]
  PIN m_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END m_in[123]
  PIN m_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END m_in[124]
  PIN m_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 456.320 4.000 456.920 ;
    END
  END m_in[125]
  PIN m_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 4.000 460.320 ;
    END
  END m_in[126]
  PIN m_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.120 4.000 463.720 ;
    END
  END m_in[127]
  PIN m_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END m_in[128]
  PIN m_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END m_in[129]
  PIN m_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END m_in[12]
  PIN m_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.000 4.000 474.600 ;
    END
  END m_in[130]
  PIN m_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 4.000 478.000 ;
    END
  END m_in[131]
  PIN m_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 4.000 55.720 ;
    END
  END m_in[13]
  PIN m_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END m_in[14]
  PIN m_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END m_in[15]
  PIN m_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END m_in[16]
  PIN m_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END m_in[17]
  PIN m_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END m_in[18]
  PIN m_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END m_in[19]
  PIN m_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END m_in[1]
  PIN m_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END m_in[20]
  PIN m_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 4.000 84.280 ;
    END
  END m_in[21]
  PIN m_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END m_in[22]
  PIN m_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END m_in[23]
  PIN m_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END m_in[24]
  PIN m_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END m_in[25]
  PIN m_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END m_in[26]
  PIN m_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END m_in[27]
  PIN m_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END m_in[28]
  PIN m_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END m_in[29]
  PIN m_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END m_in[2]
  PIN m_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END m_in[30]
  PIN m_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END m_in[31]
  PIN m_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END m_in[32]
  PIN m_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END m_in[33]
  PIN m_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END m_in[34]
  PIN m_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END m_in[35]
  PIN m_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END m_in[36]
  PIN m_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.800 4.000 141.400 ;
    END
  END m_in[37]
  PIN m_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END m_in[38]
  PIN m_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END m_in[39]
  PIN m_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END m_in[3]
  PIN m_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.680 4.000 152.280 ;
    END
  END m_in[40]
  PIN m_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END m_in[41]
  PIN m_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END m_in[42]
  PIN m_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END m_in[43]
  PIN m_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END m_in[44]
  PIN m_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 169.360 4.000 169.960 ;
    END
  END m_in[45]
  PIN m_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END m_in[46]
  PIN m_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END m_in[47]
  PIN m_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END m_in[48]
  PIN m_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END m_in[49]
  PIN m_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END m_in[4]
  PIN m_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END m_in[50]
  PIN m_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END m_in[51]
  PIN m_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END m_in[52]
  PIN m_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.920 4.000 198.520 ;
    END
  END m_in[53]
  PIN m_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END m_in[54]
  PIN m_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END m_in[55]
  PIN m_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.800 4.000 209.400 ;
    END
  END m_in[56]
  PIN m_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END m_in[57]
  PIN m_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END m_in[58]
  PIN m_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END m_in[59]
  PIN m_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END m_in[5]
  PIN m_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END m_in[60]
  PIN m_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 226.480 4.000 227.080 ;
    END
  END m_in[61]
  PIN m_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.560 4.000 231.160 ;
    END
  END m_in[62]
  PIN m_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END m_in[63]
  PIN m_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.360 4.000 237.960 ;
    END
  END m_in[64]
  PIN m_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END m_in[65]
  PIN m_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END m_in[66]
  PIN m_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END m_in[67]
  PIN m_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END m_in[68]
  PIN m_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END m_in[69]
  PIN m_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END m_in[6]
  PIN m_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END m_in[70]
  PIN m_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END m_in[71]
  PIN m_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.920 4.000 266.520 ;
    END
  END m_in[72]
  PIN m_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END m_in[73]
  PIN m_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END m_in[74]
  PIN m_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.800 4.000 277.400 ;
    END
  END m_in[75]
  PIN m_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END m_in[76]
  PIN m_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END m_in[77]
  PIN m_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.680 4.000 288.280 ;
    END
  END m_in[78]
  PIN m_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END m_in[79]
  PIN m_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END m_in[7]
  PIN m_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END m_in[80]
  PIN m_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.560 4.000 299.160 ;
    END
  END m_in[81]
  PIN m_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END m_in[82]
  PIN m_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.360 4.000 305.960 ;
    END
  END m_in[83]
  PIN m_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END m_in[84]
  PIN m_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END m_in[85]
  PIN m_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END m_in[86]
  PIN m_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END m_in[87]
  PIN m_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END m_in[88]
  PIN m_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.120 4.000 327.720 ;
    END
  END m_in[89]
  PIN m_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END m_in[8]
  PIN m_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END m_in[90]
  PIN m_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.920 4.000 334.520 ;
    END
  END m_in[91]
  PIN m_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.000 4.000 338.600 ;
    END
  END m_in[92]
  PIN m_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END m_in[93]
  PIN m_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.800 4.000 345.400 ;
    END
  END m_in[94]
  PIN m_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.880 4.000 349.480 ;
    END
  END m_in[95]
  PIN m_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END m_in[96]
  PIN m_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.680 4.000 356.280 ;
    END
  END m_in[97]
  PIN m_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END m_in[98]
  PIN m_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END m_in[99]
  PIN m_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END m_in[9]
  PIN m_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 481.480 4.000 482.080 ;
    END
  END m_out[0]
  PIN m_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END m_out[10]
  PIN m_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END m_out[11]
  PIN m_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 524.320 4.000 524.920 ;
    END
  END m_out[12]
  PIN m_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END m_out[13]
  PIN m_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.120 4.000 531.720 ;
    END
  END m_out[14]
  PIN m_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.200 4.000 535.800 ;
    END
  END m_out[15]
  PIN m_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 538.600 4.000 539.200 ;
    END
  END m_out[16]
  PIN m_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.000 4.000 542.600 ;
    END
  END m_out[17]
  PIN m_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 545.400 4.000 546.000 ;
    END
  END m_out[18]
  PIN m_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 549.480 4.000 550.080 ;
    END
  END m_out[19]
  PIN m_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.880 4.000 485.480 ;
    END
  END m_out[1]
  PIN m_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.880 4.000 553.480 ;
    END
  END m_out[20]
  PIN m_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.280 4.000 556.880 ;
    END
  END m_out[21]
  PIN m_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.680 4.000 560.280 ;
    END
  END m_out[22]
  PIN m_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.760 4.000 564.360 ;
    END
  END m_out[23]
  PIN m_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.160 4.000 567.760 ;
    END
  END m_out[24]
  PIN m_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 570.560 4.000 571.160 ;
    END
  END m_out[25]
  PIN m_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 4.000 574.560 ;
    END
  END m_out[26]
  PIN m_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END m_out[27]
  PIN m_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 581.440 4.000 582.040 ;
    END
  END m_out[28]
  PIN m_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END m_out[29]
  PIN m_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END m_out[2]
  PIN m_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.920 4.000 589.520 ;
    END
  END m_out[30]
  PIN m_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 592.320 4.000 592.920 ;
    END
  END m_out[31]
  PIN m_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.720 4.000 596.320 ;
    END
  END m_out[32]
  PIN m_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.120 4.000 599.720 ;
    END
  END m_out[33]
  PIN m_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.200 4.000 603.800 ;
    END
  END m_out[34]
  PIN m_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 606.600 4.000 607.200 ;
    END
  END m_out[35]
  PIN m_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.000 4.000 610.600 ;
    END
  END m_out[36]
  PIN m_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 613.400 4.000 614.000 ;
    END
  END m_out[37]
  PIN m_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.480 4.000 618.080 ;
    END
  END m_out[38]
  PIN m_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.880 4.000 621.480 ;
    END
  END m_out[39]
  PIN m_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.680 4.000 492.280 ;
    END
  END m_out[3]
  PIN m_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END m_out[40]
  PIN m_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 628.360 4.000 628.960 ;
    END
  END m_out[41]
  PIN m_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.760 4.000 632.360 ;
    END
  END m_out[42]
  PIN m_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.160 4.000 635.760 ;
    END
  END m_out[43]
  PIN m_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 638.560 4.000 639.160 ;
    END
  END m_out[44]
  PIN m_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END m_out[45]
  PIN m_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END m_out[46]
  PIN m_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 649.440 4.000 650.040 ;
    END
  END m_out[47]
  PIN m_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END m_out[48]
  PIN m_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.920 4.000 657.520 ;
    END
  END m_out[49]
  PIN m_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.760 4.000 496.360 ;
    END
  END m_out[4]
  PIN m_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 660.320 4.000 660.920 ;
    END
  END m_out[50]
  PIN m_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.720 4.000 664.320 ;
    END
  END m_out[51]
  PIN m_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.120 4.000 667.720 ;
    END
  END m_out[52]
  PIN m_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.200 4.000 671.800 ;
    END
  END m_out[53]
  PIN m_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 674.600 4.000 675.200 ;
    END
  END m_out[54]
  PIN m_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.000 4.000 678.600 ;
    END
  END m_out[55]
  PIN m_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 682.080 4.000 682.680 ;
    END
  END m_out[56]
  PIN m_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 685.480 4.000 686.080 ;
    END
  END m_out[57]
  PIN m_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.880 4.000 689.480 ;
    END
  END m_out[58]
  PIN m_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 692.280 4.000 692.880 ;
    END
  END m_out[59]
  PIN m_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END m_out[5]
  PIN m_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 696.360 4.000 696.960 ;
    END
  END m_out[60]
  PIN m_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.760 4.000 700.360 ;
    END
  END m_out[61]
  PIN m_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.160 4.000 703.760 ;
    END
  END m_out[62]
  PIN m_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 706.560 4.000 707.160 ;
    END
  END m_out[63]
  PIN m_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 710.640 4.000 711.240 ;
    END
  END m_out[64]
  PIN m_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END m_out[65]
  PIN m_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END m_out[66]
  PIN m_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 502.560 4.000 503.160 ;
    END
  END m_out[6]
  PIN m_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.960 4.000 506.560 ;
    END
  END m_out[7]
  PIN m_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END m_out[8]
  PIN m_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 4.000 514.040 ;
    END
  END m_out[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END rst
  PIN stall_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END stall_out
  PIN wishbone_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 716.000 2.210 720.000 ;
    END
  END wishbone_in[0]
  PIN wishbone_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 716.000 43.610 720.000 ;
    END
  END wishbone_in[10]
  PIN wishbone_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 716.000 47.750 720.000 ;
    END
  END wishbone_in[11]
  PIN wishbone_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 716.000 51.890 720.000 ;
    END
  END wishbone_in[12]
  PIN wishbone_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 716.000 56.030 720.000 ;
    END
  END wishbone_in[13]
  PIN wishbone_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 716.000 60.170 720.000 ;
    END
  END wishbone_in[14]
  PIN wishbone_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 716.000 64.310 720.000 ;
    END
  END wishbone_in[15]
  PIN wishbone_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 716.000 68.450 720.000 ;
    END
  END wishbone_in[16]
  PIN wishbone_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 716.000 72.590 720.000 ;
    END
  END wishbone_in[17]
  PIN wishbone_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 716.000 76.730 720.000 ;
    END
  END wishbone_in[18]
  PIN wishbone_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 716.000 80.870 720.000 ;
    END
  END wishbone_in[19]
  PIN wishbone_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 716.000 6.350 720.000 ;
    END
  END wishbone_in[1]
  PIN wishbone_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 716.000 85.010 720.000 ;
    END
  END wishbone_in[20]
  PIN wishbone_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 716.000 89.150 720.000 ;
    END
  END wishbone_in[21]
  PIN wishbone_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 716.000 93.750 720.000 ;
    END
  END wishbone_in[22]
  PIN wishbone_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 716.000 97.890 720.000 ;
    END
  END wishbone_in[23]
  PIN wishbone_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 716.000 102.030 720.000 ;
    END
  END wishbone_in[24]
  PIN wishbone_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 716.000 106.170 720.000 ;
    END
  END wishbone_in[25]
  PIN wishbone_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 716.000 110.310 720.000 ;
    END
  END wishbone_in[26]
  PIN wishbone_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 716.000 114.450 720.000 ;
    END
  END wishbone_in[27]
  PIN wishbone_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 716.000 118.590 720.000 ;
    END
  END wishbone_in[28]
  PIN wishbone_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 716.000 122.730 720.000 ;
    END
  END wishbone_in[29]
  PIN wishbone_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 716.000 10.490 720.000 ;
    END
  END wishbone_in[2]
  PIN wishbone_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 716.000 126.870 720.000 ;
    END
  END wishbone_in[30]
  PIN wishbone_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 716.000 131.010 720.000 ;
    END
  END wishbone_in[31]
  PIN wishbone_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 716.000 135.150 720.000 ;
    END
  END wishbone_in[32]
  PIN wishbone_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 716.000 139.290 720.000 ;
    END
  END wishbone_in[33]
  PIN wishbone_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 716.000 143.430 720.000 ;
    END
  END wishbone_in[34]
  PIN wishbone_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 716.000 147.570 720.000 ;
    END
  END wishbone_in[35]
  PIN wishbone_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 716.000 151.710 720.000 ;
    END
  END wishbone_in[36]
  PIN wishbone_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 716.000 155.850 720.000 ;
    END
  END wishbone_in[37]
  PIN wishbone_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 716.000 159.990 720.000 ;
    END
  END wishbone_in[38]
  PIN wishbone_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 716.000 164.130 720.000 ;
    END
  END wishbone_in[39]
  PIN wishbone_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 716.000 14.630 720.000 ;
    END
  END wishbone_in[3]
  PIN wishbone_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 716.000 168.270 720.000 ;
    END
  END wishbone_in[40]
  PIN wishbone_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 716.000 172.410 720.000 ;
    END
  END wishbone_in[41]
  PIN wishbone_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 716.000 176.550 720.000 ;
    END
  END wishbone_in[42]
  PIN wishbone_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 716.000 180.690 720.000 ;
    END
  END wishbone_in[43]
  PIN wishbone_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 716.000 185.290 720.000 ;
    END
  END wishbone_in[44]
  PIN wishbone_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 716.000 189.430 720.000 ;
    END
  END wishbone_in[45]
  PIN wishbone_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 716.000 193.570 720.000 ;
    END
  END wishbone_in[46]
  PIN wishbone_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 716.000 197.710 720.000 ;
    END
  END wishbone_in[47]
  PIN wishbone_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 716.000 201.850 720.000 ;
    END
  END wishbone_in[48]
  PIN wishbone_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 716.000 205.990 720.000 ;
    END
  END wishbone_in[49]
  PIN wishbone_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 716.000 18.770 720.000 ;
    END
  END wishbone_in[4]
  PIN wishbone_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 716.000 210.130 720.000 ;
    END
  END wishbone_in[50]
  PIN wishbone_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 716.000 214.270 720.000 ;
    END
  END wishbone_in[51]
  PIN wishbone_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 716.000 218.410 720.000 ;
    END
  END wishbone_in[52]
  PIN wishbone_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 716.000 222.550 720.000 ;
    END
  END wishbone_in[53]
  PIN wishbone_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 716.000 226.690 720.000 ;
    END
  END wishbone_in[54]
  PIN wishbone_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 716.000 230.830 720.000 ;
    END
  END wishbone_in[55]
  PIN wishbone_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 716.000 234.970 720.000 ;
    END
  END wishbone_in[56]
  PIN wishbone_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 716.000 239.110 720.000 ;
    END
  END wishbone_in[57]
  PIN wishbone_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 716.000 243.250 720.000 ;
    END
  END wishbone_in[58]
  PIN wishbone_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 716.000 247.390 720.000 ;
    END
  END wishbone_in[59]
  PIN wishbone_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 716.000 22.910 720.000 ;
    END
  END wishbone_in[5]
  PIN wishbone_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 716.000 251.530 720.000 ;
    END
  END wishbone_in[60]
  PIN wishbone_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 716.000 255.670 720.000 ;
    END
  END wishbone_in[61]
  PIN wishbone_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 716.000 259.810 720.000 ;
    END
  END wishbone_in[62]
  PIN wishbone_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 716.000 263.950 720.000 ;
    END
  END wishbone_in[63]
  PIN wishbone_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 716.000 268.090 720.000 ;
    END
  END wishbone_in[64]
  PIN wishbone_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 716.000 272.690 720.000 ;
    END
  END wishbone_in[65]
  PIN wishbone_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 716.000 27.050 720.000 ;
    END
  END wishbone_in[6]
  PIN wishbone_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 716.000 31.190 720.000 ;
    END
  END wishbone_in[7]
  PIN wishbone_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 716.000 35.330 720.000 ;
    END
  END wishbone_in[8]
  PIN wishbone_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 716.000 39.470 720.000 ;
    END
  END wishbone_in[9]
  PIN wishbone_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 716.000 276.830 720.000 ;
    END
  END wishbone_out[0]
  PIN wishbone_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 716.000 692.670 720.000 ;
    END
  END wishbone_out[100]
  PIN wishbone_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.530 716.000 696.810 720.000 ;
    END
  END wishbone_out[101]
  PIN wishbone_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.670 716.000 700.950 720.000 ;
    END
  END wishbone_out[102]
  PIN wishbone_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.810 716.000 705.090 720.000 ;
    END
  END wishbone_out[103]
  PIN wishbone_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.950 716.000 709.230 720.000 ;
    END
  END wishbone_out[104]
  PIN wishbone_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 716.000 713.370 720.000 ;
    END
  END wishbone_out[105]
  PIN wishbone_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.230 716.000 717.510 720.000 ;
    END
  END wishbone_out[106]
  PIN wishbone_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 716.000 318.230 720.000 ;
    END
  END wishbone_out[10]
  PIN wishbone_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 716.000 322.370 720.000 ;
    END
  END wishbone_out[11]
  PIN wishbone_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 716.000 326.510 720.000 ;
    END
  END wishbone_out[12]
  PIN wishbone_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 716.000 330.650 720.000 ;
    END
  END wishbone_out[13]
  PIN wishbone_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 716.000 334.790 720.000 ;
    END
  END wishbone_out[14]
  PIN wishbone_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 716.000 338.930 720.000 ;
    END
  END wishbone_out[15]
  PIN wishbone_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 716.000 343.070 720.000 ;
    END
  END wishbone_out[16]
  PIN wishbone_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 716.000 347.210 720.000 ;
    END
  END wishbone_out[17]
  PIN wishbone_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 716.000 351.350 720.000 ;
    END
  END wishbone_out[18]
  PIN wishbone_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 716.000 355.490 720.000 ;
    END
  END wishbone_out[19]
  PIN wishbone_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 716.000 280.970 720.000 ;
    END
  END wishbone_out[1]
  PIN wishbone_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 716.000 359.630 720.000 ;
    END
  END wishbone_out[20]
  PIN wishbone_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 716.000 364.230 720.000 ;
    END
  END wishbone_out[21]
  PIN wishbone_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 716.000 368.370 720.000 ;
    END
  END wishbone_out[22]
  PIN wishbone_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 716.000 372.510 720.000 ;
    END
  END wishbone_out[23]
  PIN wishbone_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 716.000 376.650 720.000 ;
    END
  END wishbone_out[24]
  PIN wishbone_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 716.000 380.790 720.000 ;
    END
  END wishbone_out[25]
  PIN wishbone_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 716.000 384.930 720.000 ;
    END
  END wishbone_out[26]
  PIN wishbone_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 716.000 389.070 720.000 ;
    END
  END wishbone_out[27]
  PIN wishbone_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 716.000 393.210 720.000 ;
    END
  END wishbone_out[28]
  PIN wishbone_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 716.000 397.350 720.000 ;
    END
  END wishbone_out[29]
  PIN wishbone_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 716.000 285.110 720.000 ;
    END
  END wishbone_out[2]
  PIN wishbone_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 716.000 401.490 720.000 ;
    END
  END wishbone_out[30]
  PIN wishbone_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.350 716.000 405.630 720.000 ;
    END
  END wishbone_out[31]
  PIN wishbone_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 716.000 409.770 720.000 ;
    END
  END wishbone_out[32]
  PIN wishbone_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 716.000 413.910 720.000 ;
    END
  END wishbone_out[33]
  PIN wishbone_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 716.000 418.050 720.000 ;
    END
  END wishbone_out[34]
  PIN wishbone_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 716.000 422.190 720.000 ;
    END
  END wishbone_out[35]
  PIN wishbone_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 716.000 426.330 720.000 ;
    END
  END wishbone_out[36]
  PIN wishbone_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 716.000 430.470 720.000 ;
    END
  END wishbone_out[37]
  PIN wishbone_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 716.000 434.610 720.000 ;
    END
  END wishbone_out[38]
  PIN wishbone_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 716.000 438.750 720.000 ;
    END
  END wishbone_out[39]
  PIN wishbone_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 716.000 289.250 720.000 ;
    END
  END wishbone_out[3]
  PIN wishbone_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 716.000 442.890 720.000 ;
    END
  END wishbone_out[40]
  PIN wishbone_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 716.000 447.030 720.000 ;
    END
  END wishbone_out[41]
  PIN wishbone_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 716.000 451.170 720.000 ;
    END
  END wishbone_out[42]
  PIN wishbone_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 716.000 455.770 720.000 ;
    END
  END wishbone_out[43]
  PIN wishbone_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.630 716.000 459.910 720.000 ;
    END
  END wishbone_out[44]
  PIN wishbone_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 716.000 464.050 720.000 ;
    END
  END wishbone_out[45]
  PIN wishbone_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 716.000 468.190 720.000 ;
    END
  END wishbone_out[46]
  PIN wishbone_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 716.000 472.330 720.000 ;
    END
  END wishbone_out[47]
  PIN wishbone_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 716.000 476.470 720.000 ;
    END
  END wishbone_out[48]
  PIN wishbone_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 716.000 480.610 720.000 ;
    END
  END wishbone_out[49]
  PIN wishbone_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 716.000 293.390 720.000 ;
    END
  END wishbone_out[4]
  PIN wishbone_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 716.000 484.750 720.000 ;
    END
  END wishbone_out[50]
  PIN wishbone_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 716.000 488.890 720.000 ;
    END
  END wishbone_out[51]
  PIN wishbone_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 716.000 493.030 720.000 ;
    END
  END wishbone_out[52]
  PIN wishbone_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 716.000 497.170 720.000 ;
    END
  END wishbone_out[53]
  PIN wishbone_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 716.000 501.310 720.000 ;
    END
  END wishbone_out[54]
  PIN wishbone_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 716.000 505.450 720.000 ;
    END
  END wishbone_out[55]
  PIN wishbone_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 716.000 509.590 720.000 ;
    END
  END wishbone_out[56]
  PIN wishbone_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 716.000 513.730 720.000 ;
    END
  END wishbone_out[57]
  PIN wishbone_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 716.000 517.870 720.000 ;
    END
  END wishbone_out[58]
  PIN wishbone_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 716.000 522.010 720.000 ;
    END
  END wishbone_out[59]
  PIN wishbone_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 716.000 297.530 720.000 ;
    END
  END wishbone_out[5]
  PIN wishbone_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.870 716.000 526.150 720.000 ;
    END
  END wishbone_out[60]
  PIN wishbone_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 716.000 530.290 720.000 ;
    END
  END wishbone_out[61]
  PIN wishbone_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 716.000 534.430 720.000 ;
    END
  END wishbone_out[62]
  PIN wishbone_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 716.000 538.570 720.000 ;
    END
  END wishbone_out[63]
  PIN wishbone_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 716.000 543.170 720.000 ;
    END
  END wishbone_out[64]
  PIN wishbone_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 716.000 547.310 720.000 ;
    END
  END wishbone_out[65]
  PIN wishbone_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 716.000 551.450 720.000 ;
    END
  END wishbone_out[66]
  PIN wishbone_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.310 716.000 555.590 720.000 ;
    END
  END wishbone_out[67]
  PIN wishbone_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 716.000 559.730 720.000 ;
    END
  END wishbone_out[68]
  PIN wishbone_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 716.000 563.870 720.000 ;
    END
  END wishbone_out[69]
  PIN wishbone_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 716.000 301.670 720.000 ;
    END
  END wishbone_out[6]
  PIN wishbone_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 716.000 568.010 720.000 ;
    END
  END wishbone_out[70]
  PIN wishbone_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.870 716.000 572.150 720.000 ;
    END
  END wishbone_out[71]
  PIN wishbone_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 716.000 576.290 720.000 ;
    END
  END wishbone_out[72]
  PIN wishbone_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 716.000 580.430 720.000 ;
    END
  END wishbone_out[73]
  PIN wishbone_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 716.000 584.570 720.000 ;
    END
  END wishbone_out[74]
  PIN wishbone_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.430 716.000 588.710 720.000 ;
    END
  END wishbone_out[75]
  PIN wishbone_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 716.000 592.850 720.000 ;
    END
  END wishbone_out[76]
  PIN wishbone_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.710 716.000 596.990 720.000 ;
    END
  END wishbone_out[77]
  PIN wishbone_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.850 716.000 601.130 720.000 ;
    END
  END wishbone_out[78]
  PIN wishbone_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.990 716.000 605.270 720.000 ;
    END
  END wishbone_out[79]
  PIN wishbone_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 716.000 305.810 720.000 ;
    END
  END wishbone_out[7]
  PIN wishbone_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 716.000 609.410 720.000 ;
    END
  END wishbone_out[80]
  PIN wishbone_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 716.000 613.550 720.000 ;
    END
  END wishbone_out[81]
  PIN wishbone_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 716.000 617.690 720.000 ;
    END
  END wishbone_out[82]
  PIN wishbone_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 716.000 621.830 720.000 ;
    END
  END wishbone_out[83]
  PIN wishbone_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 716.000 625.970 720.000 ;
    END
  END wishbone_out[84]
  PIN wishbone_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 716.000 630.110 720.000 ;
    END
  END wishbone_out[85]
  PIN wishbone_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 716.000 634.710 720.000 ;
    END
  END wishbone_out[86]
  PIN wishbone_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 716.000 638.850 720.000 ;
    END
  END wishbone_out[87]
  PIN wishbone_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 716.000 642.990 720.000 ;
    END
  END wishbone_out[88]
  PIN wishbone_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.850 716.000 647.130 720.000 ;
    END
  END wishbone_out[89]
  PIN wishbone_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 716.000 309.950 720.000 ;
    END
  END wishbone_out[8]
  PIN wishbone_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.990 716.000 651.270 720.000 ;
    END
  END wishbone_out[90]
  PIN wishbone_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.130 716.000 655.410 720.000 ;
    END
  END wishbone_out[91]
  PIN wishbone_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.270 716.000 659.550 720.000 ;
    END
  END wishbone_out[92]
  PIN wishbone_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 716.000 663.690 720.000 ;
    END
  END wishbone_out[93]
  PIN wishbone_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 716.000 667.830 720.000 ;
    END
  END wishbone_out[94]
  PIN wishbone_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.690 716.000 671.970 720.000 ;
    END
  END wishbone_out[95]
  PIN wishbone_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.830 716.000 676.110 720.000 ;
    END
  END wishbone_out[96]
  PIN wishbone_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 716.000 680.250 720.000 ;
    END
  END wishbone_out[97]
  PIN wishbone_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.110 716.000 684.390 720.000 ;
    END
  END wishbone_out[98]
  PIN wishbone_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 716.000 688.530 720.000 ;
    END
  END wishbone_out[99]
  PIN wishbone_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 716.000 314.090 720.000 ;
    END
  END wishbone_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 707.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 707.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 707.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 707.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 707.440 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 707.440 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 707.440 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 707.440 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 707.440 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 638.740 10.880 640.340 707.200 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 485.140 10.880 486.740 707.200 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 707.200 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 707.200 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 707.200 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 561.940 10.880 563.540 707.200 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 408.340 10.880 409.940 707.200 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 707.200 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 707.200 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 642.040 10.880 643.640 707.200 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 488.440 10.880 490.040 707.200 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.840 10.880 336.440 707.200 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 707.200 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 707.200 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 565.240 10.880 566.840 707.200 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 411.640 10.880 413.240 707.200 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 707.200 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 707.200 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 645.340 10.880 646.940 707.200 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 491.740 10.880 493.340 707.200 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 338.140 10.880 339.740 707.200 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 707.200 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 707.200 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 568.540 10.880 570.140 707.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 414.940 10.880 416.540 707.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 707.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 707.200 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 715.155 707.285 ;
      LAYER met1 ;
        RECT 1.450 6.160 717.990 710.900 ;
      LAYER met2 ;
        RECT 1.480 715.720 1.650 717.925 ;
        RECT 2.490 715.720 5.790 717.925 ;
        RECT 6.630 715.720 9.930 717.925 ;
        RECT 10.770 715.720 14.070 717.925 ;
        RECT 14.910 715.720 18.210 717.925 ;
        RECT 19.050 715.720 22.350 717.925 ;
        RECT 23.190 715.720 26.490 717.925 ;
        RECT 27.330 715.720 30.630 717.925 ;
        RECT 31.470 715.720 34.770 717.925 ;
        RECT 35.610 715.720 38.910 717.925 ;
        RECT 39.750 715.720 43.050 717.925 ;
        RECT 43.890 715.720 47.190 717.925 ;
        RECT 48.030 715.720 51.330 717.925 ;
        RECT 52.170 715.720 55.470 717.925 ;
        RECT 56.310 715.720 59.610 717.925 ;
        RECT 60.450 715.720 63.750 717.925 ;
        RECT 64.590 715.720 67.890 717.925 ;
        RECT 68.730 715.720 72.030 717.925 ;
        RECT 72.870 715.720 76.170 717.925 ;
        RECT 77.010 715.720 80.310 717.925 ;
        RECT 81.150 715.720 84.450 717.925 ;
        RECT 85.290 715.720 88.590 717.925 ;
        RECT 89.430 715.720 93.190 717.925 ;
        RECT 94.030 715.720 97.330 717.925 ;
        RECT 98.170 715.720 101.470 717.925 ;
        RECT 102.310 715.720 105.610 717.925 ;
        RECT 106.450 715.720 109.750 717.925 ;
        RECT 110.590 715.720 113.890 717.925 ;
        RECT 114.730 715.720 118.030 717.925 ;
        RECT 118.870 715.720 122.170 717.925 ;
        RECT 123.010 715.720 126.310 717.925 ;
        RECT 127.150 715.720 130.450 717.925 ;
        RECT 131.290 715.720 134.590 717.925 ;
        RECT 135.430 715.720 138.730 717.925 ;
        RECT 139.570 715.720 142.870 717.925 ;
        RECT 143.710 715.720 147.010 717.925 ;
        RECT 147.850 715.720 151.150 717.925 ;
        RECT 151.990 715.720 155.290 717.925 ;
        RECT 156.130 715.720 159.430 717.925 ;
        RECT 160.270 715.720 163.570 717.925 ;
        RECT 164.410 715.720 167.710 717.925 ;
        RECT 168.550 715.720 171.850 717.925 ;
        RECT 172.690 715.720 175.990 717.925 ;
        RECT 176.830 715.720 180.130 717.925 ;
        RECT 180.970 715.720 184.730 717.925 ;
        RECT 185.570 715.720 188.870 717.925 ;
        RECT 189.710 715.720 193.010 717.925 ;
        RECT 193.850 715.720 197.150 717.925 ;
        RECT 197.990 715.720 201.290 717.925 ;
        RECT 202.130 715.720 205.430 717.925 ;
        RECT 206.270 715.720 209.570 717.925 ;
        RECT 210.410 715.720 213.710 717.925 ;
        RECT 214.550 715.720 217.850 717.925 ;
        RECT 218.690 715.720 221.990 717.925 ;
        RECT 222.830 715.720 226.130 717.925 ;
        RECT 226.970 715.720 230.270 717.925 ;
        RECT 231.110 715.720 234.410 717.925 ;
        RECT 235.250 715.720 238.550 717.925 ;
        RECT 239.390 715.720 242.690 717.925 ;
        RECT 243.530 715.720 246.830 717.925 ;
        RECT 247.670 715.720 250.970 717.925 ;
        RECT 251.810 715.720 255.110 717.925 ;
        RECT 255.950 715.720 259.250 717.925 ;
        RECT 260.090 715.720 263.390 717.925 ;
        RECT 264.230 715.720 267.530 717.925 ;
        RECT 268.370 715.720 272.130 717.925 ;
        RECT 272.970 715.720 276.270 717.925 ;
        RECT 277.110 715.720 280.410 717.925 ;
        RECT 281.250 715.720 284.550 717.925 ;
        RECT 285.390 715.720 288.690 717.925 ;
        RECT 289.530 715.720 292.830 717.925 ;
        RECT 293.670 715.720 296.970 717.925 ;
        RECT 297.810 715.720 301.110 717.925 ;
        RECT 301.950 715.720 305.250 717.925 ;
        RECT 306.090 715.720 309.390 717.925 ;
        RECT 310.230 715.720 313.530 717.925 ;
        RECT 314.370 715.720 317.670 717.925 ;
        RECT 318.510 715.720 321.810 717.925 ;
        RECT 322.650 715.720 325.950 717.925 ;
        RECT 326.790 715.720 330.090 717.925 ;
        RECT 330.930 715.720 334.230 717.925 ;
        RECT 335.070 715.720 338.370 717.925 ;
        RECT 339.210 715.720 342.510 717.925 ;
        RECT 343.350 715.720 346.650 717.925 ;
        RECT 347.490 715.720 350.790 717.925 ;
        RECT 351.630 715.720 354.930 717.925 ;
        RECT 355.770 715.720 359.070 717.925 ;
        RECT 359.910 715.720 363.670 717.925 ;
        RECT 364.510 715.720 367.810 717.925 ;
        RECT 368.650 715.720 371.950 717.925 ;
        RECT 372.790 715.720 376.090 717.925 ;
        RECT 376.930 715.720 380.230 717.925 ;
        RECT 381.070 715.720 384.370 717.925 ;
        RECT 385.210 715.720 388.510 717.925 ;
        RECT 389.350 715.720 392.650 717.925 ;
        RECT 393.490 715.720 396.790 717.925 ;
        RECT 397.630 715.720 400.930 717.925 ;
        RECT 401.770 715.720 405.070 717.925 ;
        RECT 405.910 715.720 409.210 717.925 ;
        RECT 410.050 715.720 413.350 717.925 ;
        RECT 414.190 715.720 417.490 717.925 ;
        RECT 418.330 715.720 421.630 717.925 ;
        RECT 422.470 715.720 425.770 717.925 ;
        RECT 426.610 715.720 429.910 717.925 ;
        RECT 430.750 715.720 434.050 717.925 ;
        RECT 434.890 715.720 438.190 717.925 ;
        RECT 439.030 715.720 442.330 717.925 ;
        RECT 443.170 715.720 446.470 717.925 ;
        RECT 447.310 715.720 450.610 717.925 ;
        RECT 451.450 715.720 455.210 717.925 ;
        RECT 456.050 715.720 459.350 717.925 ;
        RECT 460.190 715.720 463.490 717.925 ;
        RECT 464.330 715.720 467.630 717.925 ;
        RECT 468.470 715.720 471.770 717.925 ;
        RECT 472.610 715.720 475.910 717.925 ;
        RECT 476.750 715.720 480.050 717.925 ;
        RECT 480.890 715.720 484.190 717.925 ;
        RECT 485.030 715.720 488.330 717.925 ;
        RECT 489.170 715.720 492.470 717.925 ;
        RECT 493.310 715.720 496.610 717.925 ;
        RECT 497.450 715.720 500.750 717.925 ;
        RECT 501.590 715.720 504.890 717.925 ;
        RECT 505.730 715.720 509.030 717.925 ;
        RECT 509.870 715.720 513.170 717.925 ;
        RECT 514.010 715.720 517.310 717.925 ;
        RECT 518.150 715.720 521.450 717.925 ;
        RECT 522.290 715.720 525.590 717.925 ;
        RECT 526.430 715.720 529.730 717.925 ;
        RECT 530.570 715.720 533.870 717.925 ;
        RECT 534.710 715.720 538.010 717.925 ;
        RECT 538.850 715.720 542.610 717.925 ;
        RECT 543.450 715.720 546.750 717.925 ;
        RECT 547.590 715.720 550.890 717.925 ;
        RECT 551.730 715.720 555.030 717.925 ;
        RECT 555.870 715.720 559.170 717.925 ;
        RECT 560.010 715.720 563.310 717.925 ;
        RECT 564.150 715.720 567.450 717.925 ;
        RECT 568.290 715.720 571.590 717.925 ;
        RECT 572.430 715.720 575.730 717.925 ;
        RECT 576.570 715.720 579.870 717.925 ;
        RECT 580.710 715.720 584.010 717.925 ;
        RECT 584.850 715.720 588.150 717.925 ;
        RECT 588.990 715.720 592.290 717.925 ;
        RECT 593.130 715.720 596.430 717.925 ;
        RECT 597.270 715.720 600.570 717.925 ;
        RECT 601.410 715.720 604.710 717.925 ;
        RECT 605.550 715.720 608.850 717.925 ;
        RECT 609.690 715.720 612.990 717.925 ;
        RECT 613.830 715.720 617.130 717.925 ;
        RECT 617.970 715.720 621.270 717.925 ;
        RECT 622.110 715.720 625.410 717.925 ;
        RECT 626.250 715.720 629.550 717.925 ;
        RECT 630.390 715.720 634.150 717.925 ;
        RECT 634.990 715.720 638.290 717.925 ;
        RECT 639.130 715.720 642.430 717.925 ;
        RECT 643.270 715.720 646.570 717.925 ;
        RECT 647.410 715.720 650.710 717.925 ;
        RECT 651.550 715.720 654.850 717.925 ;
        RECT 655.690 715.720 658.990 717.925 ;
        RECT 659.830 715.720 663.130 717.925 ;
        RECT 663.970 715.720 667.270 717.925 ;
        RECT 668.110 715.720 671.410 717.925 ;
        RECT 672.250 715.720 675.550 717.925 ;
        RECT 676.390 715.720 679.690 717.925 ;
        RECT 680.530 715.720 683.830 717.925 ;
        RECT 684.670 715.720 687.970 717.925 ;
        RECT 688.810 715.720 692.110 717.925 ;
        RECT 692.950 715.720 696.250 717.925 ;
        RECT 697.090 715.720 700.390 717.925 ;
        RECT 701.230 715.720 704.530 717.925 ;
        RECT 705.370 715.720 708.670 717.925 ;
        RECT 709.510 715.720 712.810 717.925 ;
        RECT 713.650 715.720 716.950 717.925 ;
        RECT 717.790 715.720 717.960 717.925 ;
        RECT 1.480 4.280 717.960 715.720 ;
        RECT 2.030 1.515 4.410 4.280 ;
        RECT 5.250 1.515 7.630 4.280 ;
        RECT 8.470 1.515 11.310 4.280 ;
        RECT 12.150 1.515 14.530 4.280 ;
        RECT 15.370 1.515 17.750 4.280 ;
        RECT 18.590 1.515 21.430 4.280 ;
        RECT 22.270 1.515 24.650 4.280 ;
        RECT 25.490 1.515 28.330 4.280 ;
        RECT 29.170 1.515 31.550 4.280 ;
        RECT 32.390 1.515 34.770 4.280 ;
        RECT 35.610 1.515 38.450 4.280 ;
        RECT 39.290 1.515 41.670 4.280 ;
        RECT 42.510 1.515 44.890 4.280 ;
        RECT 45.730 1.515 48.570 4.280 ;
        RECT 49.410 1.515 51.790 4.280 ;
        RECT 52.630 1.515 55.470 4.280 ;
        RECT 56.310 1.515 58.690 4.280 ;
        RECT 59.530 1.515 61.910 4.280 ;
        RECT 62.750 1.515 65.590 4.280 ;
        RECT 66.430 1.515 68.810 4.280 ;
        RECT 69.650 1.515 72.490 4.280 ;
        RECT 73.330 1.515 75.710 4.280 ;
        RECT 76.550 1.515 78.930 4.280 ;
        RECT 79.770 1.515 82.610 4.280 ;
        RECT 83.450 1.515 85.830 4.280 ;
        RECT 86.670 1.515 89.050 4.280 ;
        RECT 89.890 1.515 92.730 4.280 ;
        RECT 93.570 1.515 95.950 4.280 ;
        RECT 96.790 1.515 99.630 4.280 ;
        RECT 100.470 1.515 102.850 4.280 ;
        RECT 103.690 1.515 106.070 4.280 ;
        RECT 106.910 1.515 109.750 4.280 ;
        RECT 110.590 1.515 112.970 4.280 ;
        RECT 113.810 1.515 116.190 4.280 ;
        RECT 117.030 1.515 119.870 4.280 ;
        RECT 120.710 1.515 123.090 4.280 ;
        RECT 123.930 1.515 126.770 4.280 ;
        RECT 127.610 1.515 129.990 4.280 ;
        RECT 130.830 1.515 133.210 4.280 ;
        RECT 134.050 1.515 136.890 4.280 ;
        RECT 137.730 1.515 140.110 4.280 ;
        RECT 140.950 1.515 143.790 4.280 ;
        RECT 144.630 1.515 147.010 4.280 ;
        RECT 147.850 1.515 150.230 4.280 ;
        RECT 151.070 1.515 153.910 4.280 ;
        RECT 154.750 1.515 157.130 4.280 ;
        RECT 157.970 1.515 160.350 4.280 ;
        RECT 161.190 1.515 164.030 4.280 ;
        RECT 164.870 1.515 167.250 4.280 ;
        RECT 168.090 1.515 170.930 4.280 ;
        RECT 171.770 1.515 174.150 4.280 ;
        RECT 174.990 1.515 177.370 4.280 ;
        RECT 178.210 1.515 181.050 4.280 ;
        RECT 181.890 1.515 184.270 4.280 ;
        RECT 185.110 1.515 187.950 4.280 ;
        RECT 188.790 1.515 191.170 4.280 ;
        RECT 192.010 1.515 194.390 4.280 ;
        RECT 195.230 1.515 198.070 4.280 ;
        RECT 198.910 1.515 201.290 4.280 ;
        RECT 202.130 1.515 204.510 4.280 ;
        RECT 205.350 1.515 208.190 4.280 ;
        RECT 209.030 1.515 211.410 4.280 ;
        RECT 212.250 1.515 215.090 4.280 ;
        RECT 215.930 1.515 218.310 4.280 ;
        RECT 219.150 1.515 221.530 4.280 ;
        RECT 222.370 1.515 225.210 4.280 ;
        RECT 226.050 1.515 228.430 4.280 ;
        RECT 229.270 1.515 231.650 4.280 ;
        RECT 232.490 1.515 235.330 4.280 ;
        RECT 236.170 1.515 238.550 4.280 ;
        RECT 239.390 1.515 242.230 4.280 ;
        RECT 243.070 1.515 245.450 4.280 ;
        RECT 246.290 1.515 248.670 4.280 ;
        RECT 249.510 1.515 252.350 4.280 ;
        RECT 253.190 1.515 255.570 4.280 ;
        RECT 256.410 1.515 259.250 4.280 ;
        RECT 260.090 1.515 262.470 4.280 ;
        RECT 263.310 1.515 265.690 4.280 ;
        RECT 266.530 1.515 269.370 4.280 ;
        RECT 270.210 1.515 272.590 4.280 ;
        RECT 273.430 1.515 275.810 4.280 ;
        RECT 276.650 1.515 279.490 4.280 ;
        RECT 280.330 1.515 282.710 4.280 ;
        RECT 283.550 1.515 286.390 4.280 ;
        RECT 287.230 1.515 289.610 4.280 ;
        RECT 290.450 1.515 292.830 4.280 ;
        RECT 293.670 1.515 296.510 4.280 ;
        RECT 297.350 1.515 299.730 4.280 ;
        RECT 300.570 1.515 303.410 4.280 ;
        RECT 304.250 1.515 306.630 4.280 ;
        RECT 307.470 1.515 309.850 4.280 ;
        RECT 310.690 1.515 313.530 4.280 ;
        RECT 314.370 1.515 316.750 4.280 ;
        RECT 317.590 1.515 319.970 4.280 ;
        RECT 320.810 1.515 323.650 4.280 ;
        RECT 324.490 1.515 326.870 4.280 ;
        RECT 327.710 1.515 330.550 4.280 ;
        RECT 331.390 1.515 333.770 4.280 ;
        RECT 334.610 1.515 336.990 4.280 ;
        RECT 337.830 1.515 340.670 4.280 ;
        RECT 341.510 1.515 343.890 4.280 ;
        RECT 344.730 1.515 347.110 4.280 ;
        RECT 347.950 1.515 350.790 4.280 ;
        RECT 351.630 1.515 354.010 4.280 ;
        RECT 354.850 1.515 357.690 4.280 ;
        RECT 358.530 1.515 360.910 4.280 ;
        RECT 361.750 1.515 364.130 4.280 ;
        RECT 364.970 1.515 367.810 4.280 ;
        RECT 368.650 1.515 371.030 4.280 ;
        RECT 371.870 1.515 374.710 4.280 ;
        RECT 375.550 1.515 377.930 4.280 ;
        RECT 378.770 1.515 381.150 4.280 ;
        RECT 381.990 1.515 384.830 4.280 ;
        RECT 385.670 1.515 388.050 4.280 ;
        RECT 388.890 1.515 391.270 4.280 ;
        RECT 392.110 1.515 394.950 4.280 ;
        RECT 395.790 1.515 398.170 4.280 ;
        RECT 399.010 1.515 401.850 4.280 ;
        RECT 402.690 1.515 405.070 4.280 ;
        RECT 405.910 1.515 408.290 4.280 ;
        RECT 409.130 1.515 411.970 4.280 ;
        RECT 412.810 1.515 415.190 4.280 ;
        RECT 416.030 1.515 418.410 4.280 ;
        RECT 419.250 1.515 422.090 4.280 ;
        RECT 422.930 1.515 425.310 4.280 ;
        RECT 426.150 1.515 428.990 4.280 ;
        RECT 429.830 1.515 432.210 4.280 ;
        RECT 433.050 1.515 435.430 4.280 ;
        RECT 436.270 1.515 439.110 4.280 ;
        RECT 439.950 1.515 442.330 4.280 ;
        RECT 443.170 1.515 446.010 4.280 ;
        RECT 446.850 1.515 449.230 4.280 ;
        RECT 450.070 1.515 452.450 4.280 ;
        RECT 453.290 1.515 456.130 4.280 ;
        RECT 456.970 1.515 459.350 4.280 ;
        RECT 460.190 1.515 462.570 4.280 ;
        RECT 463.410 1.515 466.250 4.280 ;
        RECT 467.090 1.515 469.470 4.280 ;
        RECT 470.310 1.515 473.150 4.280 ;
        RECT 473.990 1.515 476.370 4.280 ;
        RECT 477.210 1.515 479.590 4.280 ;
        RECT 480.430 1.515 483.270 4.280 ;
        RECT 484.110 1.515 486.490 4.280 ;
        RECT 487.330 1.515 490.170 4.280 ;
        RECT 491.010 1.515 493.390 4.280 ;
        RECT 494.230 1.515 496.610 4.280 ;
        RECT 497.450 1.515 500.290 4.280 ;
        RECT 501.130 1.515 503.510 4.280 ;
        RECT 504.350 1.515 506.730 4.280 ;
        RECT 507.570 1.515 510.410 4.280 ;
        RECT 511.250 1.515 513.630 4.280 ;
        RECT 514.470 1.515 517.310 4.280 ;
        RECT 518.150 1.515 520.530 4.280 ;
        RECT 521.370 1.515 523.750 4.280 ;
        RECT 524.590 1.515 527.430 4.280 ;
        RECT 528.270 1.515 530.650 4.280 ;
        RECT 531.490 1.515 533.870 4.280 ;
        RECT 534.710 1.515 537.550 4.280 ;
        RECT 538.390 1.515 540.770 4.280 ;
        RECT 541.610 1.515 544.450 4.280 ;
        RECT 545.290 1.515 547.670 4.280 ;
        RECT 548.510 1.515 550.890 4.280 ;
        RECT 551.730 1.515 554.570 4.280 ;
        RECT 555.410 1.515 557.790 4.280 ;
        RECT 558.630 1.515 561.470 4.280 ;
        RECT 562.310 1.515 564.690 4.280 ;
        RECT 565.530 1.515 567.910 4.280 ;
        RECT 568.750 1.515 571.590 4.280 ;
        RECT 572.430 1.515 574.810 4.280 ;
        RECT 575.650 1.515 578.030 4.280 ;
        RECT 578.870 1.515 581.710 4.280 ;
        RECT 582.550 1.515 584.930 4.280 ;
        RECT 585.770 1.515 588.610 4.280 ;
        RECT 589.450 1.515 591.830 4.280 ;
        RECT 592.670 1.515 595.050 4.280 ;
        RECT 595.890 1.515 598.730 4.280 ;
        RECT 599.570 1.515 601.950 4.280 ;
        RECT 602.790 1.515 605.630 4.280 ;
        RECT 606.470 1.515 608.850 4.280 ;
        RECT 609.690 1.515 612.070 4.280 ;
        RECT 612.910 1.515 615.750 4.280 ;
        RECT 616.590 1.515 618.970 4.280 ;
        RECT 619.810 1.515 622.190 4.280 ;
        RECT 623.030 1.515 625.870 4.280 ;
        RECT 626.710 1.515 629.090 4.280 ;
        RECT 629.930 1.515 632.770 4.280 ;
        RECT 633.610 1.515 635.990 4.280 ;
        RECT 636.830 1.515 639.210 4.280 ;
        RECT 640.050 1.515 642.890 4.280 ;
        RECT 643.730 1.515 646.110 4.280 ;
        RECT 646.950 1.515 649.330 4.280 ;
        RECT 650.170 1.515 653.010 4.280 ;
        RECT 653.850 1.515 656.230 4.280 ;
        RECT 657.070 1.515 659.910 4.280 ;
        RECT 660.750 1.515 663.130 4.280 ;
        RECT 663.970 1.515 666.350 4.280 ;
        RECT 667.190 1.515 670.030 4.280 ;
        RECT 670.870 1.515 673.250 4.280 ;
        RECT 674.090 1.515 676.930 4.280 ;
        RECT 677.770 1.515 680.150 4.280 ;
        RECT 680.990 1.515 683.370 4.280 ;
        RECT 684.210 1.515 687.050 4.280 ;
        RECT 687.890 1.515 690.270 4.280 ;
        RECT 691.110 1.515 693.490 4.280 ;
        RECT 694.330 1.515 697.170 4.280 ;
        RECT 698.010 1.515 700.390 4.280 ;
        RECT 701.230 1.515 704.070 4.280 ;
        RECT 704.910 1.515 707.290 4.280 ;
        RECT 708.130 1.515 710.510 4.280 ;
        RECT 711.350 1.515 714.190 4.280 ;
        RECT 715.030 1.515 717.410 4.280 ;
      LAYER met3 ;
        RECT 4.400 717.040 714.775 717.905 ;
        RECT 3.990 715.040 714.775 717.040 ;
        RECT 4.400 713.640 714.775 715.040 ;
        RECT 3.990 711.640 714.775 713.640 ;
        RECT 4.400 710.240 714.775 711.640 ;
        RECT 3.990 707.560 714.775 710.240 ;
        RECT 4.400 706.160 714.775 707.560 ;
        RECT 3.990 704.160 714.775 706.160 ;
        RECT 4.400 702.760 714.775 704.160 ;
        RECT 3.990 700.760 714.775 702.760 ;
        RECT 4.400 699.360 714.775 700.760 ;
        RECT 3.990 697.360 714.775 699.360 ;
        RECT 4.400 695.960 714.775 697.360 ;
        RECT 3.990 693.280 714.775 695.960 ;
        RECT 4.400 691.880 714.775 693.280 ;
        RECT 3.990 689.880 714.775 691.880 ;
        RECT 4.400 688.480 714.775 689.880 ;
        RECT 3.990 686.480 714.775 688.480 ;
        RECT 4.400 685.080 714.775 686.480 ;
        RECT 3.990 683.080 714.775 685.080 ;
        RECT 4.400 681.680 714.775 683.080 ;
        RECT 3.990 679.000 714.775 681.680 ;
        RECT 4.400 677.600 714.775 679.000 ;
        RECT 3.990 675.600 714.775 677.600 ;
        RECT 4.400 674.200 714.775 675.600 ;
        RECT 3.990 672.200 714.775 674.200 ;
        RECT 4.400 670.800 714.775 672.200 ;
        RECT 3.990 668.120 714.775 670.800 ;
        RECT 4.400 666.720 714.775 668.120 ;
        RECT 3.990 664.720 714.775 666.720 ;
        RECT 4.400 663.320 714.775 664.720 ;
        RECT 3.990 661.320 714.775 663.320 ;
        RECT 4.400 659.920 714.775 661.320 ;
        RECT 3.990 657.920 714.775 659.920 ;
        RECT 4.400 656.520 714.775 657.920 ;
        RECT 3.990 653.840 714.775 656.520 ;
        RECT 4.400 652.440 714.775 653.840 ;
        RECT 3.990 650.440 714.775 652.440 ;
        RECT 4.400 649.040 714.775 650.440 ;
        RECT 3.990 647.040 714.775 649.040 ;
        RECT 4.400 645.640 714.775 647.040 ;
        RECT 3.990 643.640 714.775 645.640 ;
        RECT 4.400 642.240 714.775 643.640 ;
        RECT 3.990 639.560 714.775 642.240 ;
        RECT 4.400 638.160 714.775 639.560 ;
        RECT 3.990 636.160 714.775 638.160 ;
        RECT 4.400 634.760 714.775 636.160 ;
        RECT 3.990 632.760 714.775 634.760 ;
        RECT 4.400 631.360 714.775 632.760 ;
        RECT 3.990 629.360 714.775 631.360 ;
        RECT 4.400 627.960 714.775 629.360 ;
        RECT 3.990 625.280 714.775 627.960 ;
        RECT 4.400 623.880 714.775 625.280 ;
        RECT 3.990 621.880 714.775 623.880 ;
        RECT 4.400 620.480 714.775 621.880 ;
        RECT 3.990 618.480 714.775 620.480 ;
        RECT 4.400 617.080 714.775 618.480 ;
        RECT 3.990 614.400 714.775 617.080 ;
        RECT 4.400 613.000 714.775 614.400 ;
        RECT 3.990 611.000 714.775 613.000 ;
        RECT 4.400 609.600 714.775 611.000 ;
        RECT 3.990 607.600 714.775 609.600 ;
        RECT 4.400 606.200 714.775 607.600 ;
        RECT 3.990 604.200 714.775 606.200 ;
        RECT 4.400 602.800 714.775 604.200 ;
        RECT 3.990 600.120 714.775 602.800 ;
        RECT 4.400 598.720 714.775 600.120 ;
        RECT 3.990 596.720 714.775 598.720 ;
        RECT 4.400 595.320 714.775 596.720 ;
        RECT 3.990 593.320 714.775 595.320 ;
        RECT 4.400 591.920 714.775 593.320 ;
        RECT 3.990 589.920 714.775 591.920 ;
        RECT 4.400 588.520 714.775 589.920 ;
        RECT 3.990 585.840 714.775 588.520 ;
        RECT 4.400 584.440 714.775 585.840 ;
        RECT 3.990 582.440 714.775 584.440 ;
        RECT 4.400 581.040 714.775 582.440 ;
        RECT 3.990 579.040 714.775 581.040 ;
        RECT 4.400 577.640 714.775 579.040 ;
        RECT 3.990 574.960 714.775 577.640 ;
        RECT 4.400 573.560 714.775 574.960 ;
        RECT 3.990 571.560 714.775 573.560 ;
        RECT 4.400 570.160 714.775 571.560 ;
        RECT 3.990 568.160 714.775 570.160 ;
        RECT 4.400 566.760 714.775 568.160 ;
        RECT 3.990 564.760 714.775 566.760 ;
        RECT 4.400 563.360 714.775 564.760 ;
        RECT 3.990 560.680 714.775 563.360 ;
        RECT 4.400 559.280 714.775 560.680 ;
        RECT 3.990 557.280 714.775 559.280 ;
        RECT 4.400 555.880 714.775 557.280 ;
        RECT 3.990 553.880 714.775 555.880 ;
        RECT 4.400 552.480 714.775 553.880 ;
        RECT 3.990 550.480 714.775 552.480 ;
        RECT 4.400 549.080 714.775 550.480 ;
        RECT 3.990 546.400 714.775 549.080 ;
        RECT 4.400 545.000 714.775 546.400 ;
        RECT 3.990 543.000 714.775 545.000 ;
        RECT 4.400 541.600 714.775 543.000 ;
        RECT 3.990 539.600 714.775 541.600 ;
        RECT 4.400 538.200 714.775 539.600 ;
        RECT 3.990 536.200 714.775 538.200 ;
        RECT 4.400 534.800 714.775 536.200 ;
        RECT 3.990 532.120 714.775 534.800 ;
        RECT 4.400 530.720 714.775 532.120 ;
        RECT 3.990 528.720 714.775 530.720 ;
        RECT 4.400 527.320 714.775 528.720 ;
        RECT 3.990 525.320 714.775 527.320 ;
        RECT 4.400 523.920 714.775 525.320 ;
        RECT 3.990 521.240 714.775 523.920 ;
        RECT 4.400 519.840 714.775 521.240 ;
        RECT 3.990 517.840 714.775 519.840 ;
        RECT 4.400 516.440 714.775 517.840 ;
        RECT 3.990 514.440 714.775 516.440 ;
        RECT 4.400 513.040 714.775 514.440 ;
        RECT 3.990 511.040 714.775 513.040 ;
        RECT 4.400 509.640 714.775 511.040 ;
        RECT 3.990 506.960 714.775 509.640 ;
        RECT 4.400 505.560 714.775 506.960 ;
        RECT 3.990 503.560 714.775 505.560 ;
        RECT 4.400 502.160 714.775 503.560 ;
        RECT 3.990 500.160 714.775 502.160 ;
        RECT 4.400 498.760 714.775 500.160 ;
        RECT 3.990 496.760 714.775 498.760 ;
        RECT 4.400 495.360 714.775 496.760 ;
        RECT 3.990 492.680 714.775 495.360 ;
        RECT 4.400 491.280 714.775 492.680 ;
        RECT 3.990 489.280 714.775 491.280 ;
        RECT 4.400 487.880 714.775 489.280 ;
        RECT 3.990 485.880 714.775 487.880 ;
        RECT 4.400 484.480 714.775 485.880 ;
        RECT 3.990 482.480 714.775 484.480 ;
        RECT 4.400 481.080 714.775 482.480 ;
        RECT 3.990 478.400 714.775 481.080 ;
        RECT 4.400 477.000 714.775 478.400 ;
        RECT 3.990 475.000 714.775 477.000 ;
        RECT 4.400 473.600 714.775 475.000 ;
        RECT 3.990 471.600 714.775 473.600 ;
        RECT 4.400 470.200 714.775 471.600 ;
        RECT 3.990 467.520 714.775 470.200 ;
        RECT 4.400 466.120 714.775 467.520 ;
        RECT 3.990 464.120 714.775 466.120 ;
        RECT 4.400 462.720 714.775 464.120 ;
        RECT 3.990 460.720 714.775 462.720 ;
        RECT 4.400 459.320 714.775 460.720 ;
        RECT 3.990 457.320 714.775 459.320 ;
        RECT 4.400 455.920 714.775 457.320 ;
        RECT 3.990 453.240 714.775 455.920 ;
        RECT 4.400 451.840 714.775 453.240 ;
        RECT 3.990 449.840 714.775 451.840 ;
        RECT 4.400 448.440 714.775 449.840 ;
        RECT 3.990 446.440 714.775 448.440 ;
        RECT 4.400 445.040 714.775 446.440 ;
        RECT 3.990 443.040 714.775 445.040 ;
        RECT 4.400 441.640 714.775 443.040 ;
        RECT 3.990 438.960 714.775 441.640 ;
        RECT 4.400 437.560 714.775 438.960 ;
        RECT 3.990 435.560 714.775 437.560 ;
        RECT 4.400 434.160 714.775 435.560 ;
        RECT 3.990 432.160 714.775 434.160 ;
        RECT 4.400 430.760 714.775 432.160 ;
        RECT 3.990 428.080 714.775 430.760 ;
        RECT 4.400 426.680 714.775 428.080 ;
        RECT 3.990 424.680 714.775 426.680 ;
        RECT 4.400 423.280 714.775 424.680 ;
        RECT 3.990 421.280 714.775 423.280 ;
        RECT 4.400 419.880 714.775 421.280 ;
        RECT 3.990 417.880 714.775 419.880 ;
        RECT 4.400 416.480 714.775 417.880 ;
        RECT 3.990 413.800 714.775 416.480 ;
        RECT 4.400 412.400 714.775 413.800 ;
        RECT 3.990 410.400 714.775 412.400 ;
        RECT 4.400 409.000 714.775 410.400 ;
        RECT 3.990 407.000 714.775 409.000 ;
        RECT 4.400 405.600 714.775 407.000 ;
        RECT 3.990 403.600 714.775 405.600 ;
        RECT 4.400 402.200 714.775 403.600 ;
        RECT 3.990 399.520 714.775 402.200 ;
        RECT 4.400 398.120 714.775 399.520 ;
        RECT 3.990 396.120 714.775 398.120 ;
        RECT 4.400 394.720 714.775 396.120 ;
        RECT 3.990 392.720 714.775 394.720 ;
        RECT 4.400 391.320 714.775 392.720 ;
        RECT 3.990 389.320 714.775 391.320 ;
        RECT 4.400 387.920 714.775 389.320 ;
        RECT 3.990 385.240 714.775 387.920 ;
        RECT 4.400 383.840 714.775 385.240 ;
        RECT 3.990 381.840 714.775 383.840 ;
        RECT 4.400 380.440 714.775 381.840 ;
        RECT 3.990 378.440 714.775 380.440 ;
        RECT 4.400 377.040 714.775 378.440 ;
        RECT 3.990 374.360 714.775 377.040 ;
        RECT 4.400 372.960 714.775 374.360 ;
        RECT 3.990 370.960 714.775 372.960 ;
        RECT 4.400 369.560 714.775 370.960 ;
        RECT 3.990 367.560 714.775 369.560 ;
        RECT 4.400 366.160 714.775 367.560 ;
        RECT 3.990 364.160 714.775 366.160 ;
        RECT 4.400 362.760 714.775 364.160 ;
        RECT 3.990 360.080 714.775 362.760 ;
        RECT 4.400 358.680 714.775 360.080 ;
        RECT 3.990 356.680 714.775 358.680 ;
        RECT 4.400 355.280 714.775 356.680 ;
        RECT 3.990 353.280 714.775 355.280 ;
        RECT 4.400 351.880 714.775 353.280 ;
        RECT 3.990 349.880 714.775 351.880 ;
        RECT 4.400 348.480 714.775 349.880 ;
        RECT 3.990 345.800 714.775 348.480 ;
        RECT 4.400 344.400 714.775 345.800 ;
        RECT 3.990 342.400 714.775 344.400 ;
        RECT 4.400 341.000 714.775 342.400 ;
        RECT 3.990 339.000 714.775 341.000 ;
        RECT 4.400 337.600 714.775 339.000 ;
        RECT 3.990 334.920 714.775 337.600 ;
        RECT 4.400 333.520 714.775 334.920 ;
        RECT 3.990 331.520 714.775 333.520 ;
        RECT 4.400 330.120 714.775 331.520 ;
        RECT 3.990 328.120 714.775 330.120 ;
        RECT 4.400 326.720 714.775 328.120 ;
        RECT 3.990 324.720 714.775 326.720 ;
        RECT 4.400 323.320 714.775 324.720 ;
        RECT 3.990 320.640 714.775 323.320 ;
        RECT 4.400 319.240 714.775 320.640 ;
        RECT 3.990 317.240 714.775 319.240 ;
        RECT 4.400 315.840 714.775 317.240 ;
        RECT 3.990 313.840 714.775 315.840 ;
        RECT 4.400 312.440 714.775 313.840 ;
        RECT 3.990 310.440 714.775 312.440 ;
        RECT 4.400 309.040 714.775 310.440 ;
        RECT 3.990 306.360 714.775 309.040 ;
        RECT 4.400 304.960 714.775 306.360 ;
        RECT 3.990 302.960 714.775 304.960 ;
        RECT 4.400 301.560 714.775 302.960 ;
        RECT 3.990 299.560 714.775 301.560 ;
        RECT 4.400 298.160 714.775 299.560 ;
        RECT 3.990 296.160 714.775 298.160 ;
        RECT 4.400 294.760 714.775 296.160 ;
        RECT 3.990 292.080 714.775 294.760 ;
        RECT 4.400 290.680 714.775 292.080 ;
        RECT 3.990 288.680 714.775 290.680 ;
        RECT 4.400 287.280 714.775 288.680 ;
        RECT 3.990 285.280 714.775 287.280 ;
        RECT 4.400 283.880 714.775 285.280 ;
        RECT 3.990 281.200 714.775 283.880 ;
        RECT 4.400 279.800 714.775 281.200 ;
        RECT 3.990 277.800 714.775 279.800 ;
        RECT 4.400 276.400 714.775 277.800 ;
        RECT 3.990 274.400 714.775 276.400 ;
        RECT 4.400 273.000 714.775 274.400 ;
        RECT 3.990 271.000 714.775 273.000 ;
        RECT 4.400 269.600 714.775 271.000 ;
        RECT 3.990 266.920 714.775 269.600 ;
        RECT 4.400 265.520 714.775 266.920 ;
        RECT 3.990 263.520 714.775 265.520 ;
        RECT 4.400 262.120 714.775 263.520 ;
        RECT 3.990 260.120 714.775 262.120 ;
        RECT 4.400 258.720 714.775 260.120 ;
        RECT 3.990 256.720 714.775 258.720 ;
        RECT 4.400 255.320 714.775 256.720 ;
        RECT 3.990 252.640 714.775 255.320 ;
        RECT 4.400 251.240 714.775 252.640 ;
        RECT 3.990 249.240 714.775 251.240 ;
        RECT 4.400 247.840 714.775 249.240 ;
        RECT 3.990 245.840 714.775 247.840 ;
        RECT 4.400 244.440 714.775 245.840 ;
        RECT 3.990 242.440 714.775 244.440 ;
        RECT 4.400 241.040 714.775 242.440 ;
        RECT 3.990 238.360 714.775 241.040 ;
        RECT 4.400 236.960 714.775 238.360 ;
        RECT 3.990 234.960 714.775 236.960 ;
        RECT 4.400 233.560 714.775 234.960 ;
        RECT 3.990 231.560 714.775 233.560 ;
        RECT 4.400 230.160 714.775 231.560 ;
        RECT 3.990 227.480 714.775 230.160 ;
        RECT 4.400 226.080 714.775 227.480 ;
        RECT 3.990 224.080 714.775 226.080 ;
        RECT 4.400 222.680 714.775 224.080 ;
        RECT 3.990 220.680 714.775 222.680 ;
        RECT 4.400 219.280 714.775 220.680 ;
        RECT 3.990 217.280 714.775 219.280 ;
        RECT 4.400 215.880 714.775 217.280 ;
        RECT 3.990 213.200 714.775 215.880 ;
        RECT 4.400 211.800 714.775 213.200 ;
        RECT 3.990 209.800 714.775 211.800 ;
        RECT 4.400 208.400 714.775 209.800 ;
        RECT 3.990 206.400 714.775 208.400 ;
        RECT 4.400 205.000 714.775 206.400 ;
        RECT 3.990 203.000 714.775 205.000 ;
        RECT 4.400 201.600 714.775 203.000 ;
        RECT 3.990 198.920 714.775 201.600 ;
        RECT 4.400 197.520 714.775 198.920 ;
        RECT 3.990 195.520 714.775 197.520 ;
        RECT 4.400 194.120 714.775 195.520 ;
        RECT 3.990 192.120 714.775 194.120 ;
        RECT 4.400 190.720 714.775 192.120 ;
        RECT 3.990 188.040 714.775 190.720 ;
        RECT 4.400 186.640 714.775 188.040 ;
        RECT 3.990 184.640 714.775 186.640 ;
        RECT 4.400 183.240 714.775 184.640 ;
        RECT 3.990 181.240 714.775 183.240 ;
        RECT 4.400 179.840 714.775 181.240 ;
        RECT 3.990 177.840 714.775 179.840 ;
        RECT 4.400 176.440 714.775 177.840 ;
        RECT 3.990 173.760 714.775 176.440 ;
        RECT 4.400 172.360 714.775 173.760 ;
        RECT 3.990 170.360 714.775 172.360 ;
        RECT 4.400 168.960 714.775 170.360 ;
        RECT 3.990 166.960 714.775 168.960 ;
        RECT 4.400 165.560 714.775 166.960 ;
        RECT 3.990 163.560 714.775 165.560 ;
        RECT 4.400 162.160 714.775 163.560 ;
        RECT 3.990 159.480 714.775 162.160 ;
        RECT 4.400 158.080 714.775 159.480 ;
        RECT 3.990 156.080 714.775 158.080 ;
        RECT 4.400 154.680 714.775 156.080 ;
        RECT 3.990 152.680 714.775 154.680 ;
        RECT 4.400 151.280 714.775 152.680 ;
        RECT 3.990 149.280 714.775 151.280 ;
        RECT 4.400 147.880 714.775 149.280 ;
        RECT 3.990 145.200 714.775 147.880 ;
        RECT 4.400 143.800 714.775 145.200 ;
        RECT 3.990 141.800 714.775 143.800 ;
        RECT 4.400 140.400 714.775 141.800 ;
        RECT 3.990 138.400 714.775 140.400 ;
        RECT 4.400 137.000 714.775 138.400 ;
        RECT 3.990 134.320 714.775 137.000 ;
        RECT 4.400 132.920 714.775 134.320 ;
        RECT 3.990 130.920 714.775 132.920 ;
        RECT 4.400 129.520 714.775 130.920 ;
        RECT 3.990 127.520 714.775 129.520 ;
        RECT 4.400 126.120 714.775 127.520 ;
        RECT 3.990 124.120 714.775 126.120 ;
        RECT 4.400 122.720 714.775 124.120 ;
        RECT 3.990 120.040 714.775 122.720 ;
        RECT 4.400 118.640 714.775 120.040 ;
        RECT 3.990 116.640 714.775 118.640 ;
        RECT 4.400 115.240 714.775 116.640 ;
        RECT 3.990 113.240 714.775 115.240 ;
        RECT 4.400 111.840 714.775 113.240 ;
        RECT 3.990 109.840 714.775 111.840 ;
        RECT 4.400 108.440 714.775 109.840 ;
        RECT 3.990 105.760 714.775 108.440 ;
        RECT 4.400 104.360 714.775 105.760 ;
        RECT 3.990 102.360 714.775 104.360 ;
        RECT 4.400 100.960 714.775 102.360 ;
        RECT 3.990 98.960 714.775 100.960 ;
        RECT 4.400 97.560 714.775 98.960 ;
        RECT 3.990 94.880 714.775 97.560 ;
        RECT 4.400 93.480 714.775 94.880 ;
        RECT 3.990 91.480 714.775 93.480 ;
        RECT 4.400 90.080 714.775 91.480 ;
        RECT 3.990 88.080 714.775 90.080 ;
        RECT 4.400 86.680 714.775 88.080 ;
        RECT 3.990 84.680 714.775 86.680 ;
        RECT 4.400 83.280 714.775 84.680 ;
        RECT 3.990 80.600 714.775 83.280 ;
        RECT 4.400 79.200 714.775 80.600 ;
        RECT 3.990 77.200 714.775 79.200 ;
        RECT 4.400 75.800 714.775 77.200 ;
        RECT 3.990 73.800 714.775 75.800 ;
        RECT 4.400 72.400 714.775 73.800 ;
        RECT 3.990 70.400 714.775 72.400 ;
        RECT 4.400 69.000 714.775 70.400 ;
        RECT 3.990 66.320 714.775 69.000 ;
        RECT 4.400 64.920 714.775 66.320 ;
        RECT 3.990 62.920 714.775 64.920 ;
        RECT 4.400 61.520 714.775 62.920 ;
        RECT 3.990 59.520 714.775 61.520 ;
        RECT 4.400 58.120 714.775 59.520 ;
        RECT 3.990 56.120 714.775 58.120 ;
        RECT 4.400 54.720 714.775 56.120 ;
        RECT 3.990 52.040 714.775 54.720 ;
        RECT 4.400 50.640 714.775 52.040 ;
        RECT 3.990 48.640 714.775 50.640 ;
        RECT 4.400 47.240 714.775 48.640 ;
        RECT 3.990 45.240 714.775 47.240 ;
        RECT 4.400 43.840 714.775 45.240 ;
        RECT 3.990 41.160 714.775 43.840 ;
        RECT 4.400 39.760 714.775 41.160 ;
        RECT 3.990 37.760 714.775 39.760 ;
        RECT 4.400 36.360 714.775 37.760 ;
        RECT 3.990 34.360 714.775 36.360 ;
        RECT 4.400 32.960 714.775 34.360 ;
        RECT 3.990 30.960 714.775 32.960 ;
        RECT 4.400 29.560 714.775 30.960 ;
        RECT 3.990 26.880 714.775 29.560 ;
        RECT 4.400 25.480 714.775 26.880 ;
        RECT 3.990 23.480 714.775 25.480 ;
        RECT 4.400 22.080 714.775 23.480 ;
        RECT 3.990 20.080 714.775 22.080 ;
        RECT 4.400 18.680 714.775 20.080 ;
        RECT 3.990 16.680 714.775 18.680 ;
        RECT 4.400 15.280 714.775 16.680 ;
        RECT 3.990 12.600 714.775 15.280 ;
        RECT 4.400 11.200 714.775 12.600 ;
        RECT 3.990 9.200 714.775 11.200 ;
        RECT 4.400 7.800 714.775 9.200 ;
        RECT 3.990 5.800 714.775 7.800 ;
        RECT 4.400 4.400 714.775 5.800 ;
        RECT 3.990 2.400 714.775 4.400 ;
        RECT 4.400 1.535 714.775 2.400 ;
      LAYER met4 ;
        RECT 37.095 707.840 678.665 715.865 ;
        RECT 37.095 13.095 97.440 707.840 ;
        RECT 99.840 707.600 174.240 707.840 ;
        RECT 99.840 13.095 100.740 707.600 ;
        RECT 103.140 13.095 104.040 707.600 ;
        RECT 106.440 13.095 107.340 707.600 ;
        RECT 109.740 13.095 174.240 707.600 ;
        RECT 176.640 707.600 251.040 707.840 ;
        RECT 176.640 13.095 177.540 707.600 ;
        RECT 179.940 13.095 180.840 707.600 ;
        RECT 183.240 13.095 184.140 707.600 ;
        RECT 186.540 13.095 251.040 707.600 ;
        RECT 253.440 707.600 327.840 707.840 ;
        RECT 253.440 13.095 254.340 707.600 ;
        RECT 256.740 13.095 257.640 707.600 ;
        RECT 260.040 13.095 260.940 707.600 ;
        RECT 263.340 13.095 327.840 707.600 ;
        RECT 330.240 707.600 404.640 707.840 ;
        RECT 330.240 13.095 331.140 707.600 ;
        RECT 333.540 13.095 334.440 707.600 ;
        RECT 336.840 13.095 337.740 707.600 ;
        RECT 340.140 13.095 404.640 707.600 ;
        RECT 407.040 707.600 481.440 707.840 ;
        RECT 407.040 13.095 407.940 707.600 ;
        RECT 410.340 13.095 411.240 707.600 ;
        RECT 413.640 13.095 414.540 707.600 ;
        RECT 416.940 13.095 481.440 707.600 ;
        RECT 483.840 707.600 558.240 707.840 ;
        RECT 483.840 13.095 484.740 707.600 ;
        RECT 487.140 13.095 488.040 707.600 ;
        RECT 490.440 13.095 491.340 707.600 ;
        RECT 493.740 13.095 558.240 707.600 ;
        RECT 560.640 707.600 635.040 707.840 ;
        RECT 560.640 13.095 561.540 707.600 ;
        RECT 563.940 13.095 564.840 707.600 ;
        RECT 567.240 13.095 568.140 707.600 ;
        RECT 570.540 13.095 635.040 707.600 ;
        RECT 637.440 707.600 678.665 707.840 ;
        RECT 637.440 13.095 638.340 707.600 ;
        RECT 640.740 13.095 641.640 707.600 ;
        RECT 644.040 13.095 644.940 707.600 ;
        RECT 647.340 13.095 678.665 707.600 ;
  END
END dcache
END LIBRARY

